************************************************************************
* auCdl Netlist:
* 
* Library Name:  SRAM_ChargePulsation
* Top Cell Name: SRAMCIMfinal
* View Name:     schematic
* Netlisted on:  Aug 21 21:42:47 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

.lib '/data/home/chentingran/PDK/SPDK55LL_ULP_09121825_OA_CDS_V1.15_0/smic55ll_ulp_09121825_oa_cds_v1.15_0/models/hspice/l0055ll_v1p15.lib' TT
.lib '/data/home/chentingran/PDK/SPDK55LL_ULP_09121825_OA_CDS_V1.15_0/smic55ll_ulp_09121825_oa_cds_v1.15_0/models/hspice/l0055ll_v1p15.lib' RES_TT
.lib '/data/home/chentingran/PDK/SPDK55LL_ULP_09121825_OA_CDS_V1.15_0/smic55ll_ulp_09121825_oa_cds_v1.15_0/models/hspice/l0055ll_v1p15.lib' MOM_TT
.options MACMOD=1


************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    cell_SRAM
* View Name:    schematic
************************************************************************

.SUBCKT cell_SRAM BL Q QN SL VDD VSS WL
*.PININFO WL:I Q:O QN:O BL:B SL:B VDD:B VSS:B
XPM0 QN Q VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM1 Q QN VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XNM5 Q QN VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM4 QN Q VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM3 Q WL SL VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM2 BL WL QN VSS n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    cell_PIM
* View Name:    schematic
************************************************************************

.SUBCKT cell_PIM bl cbl in1 in2 sl vdd vss wl
*.PININFO bl:I in1:I in2:I sl:I wl:I cbl:B vdd:B vss:B
XI0 bl q qn sl vdd vss wl / cell_SRAM
XM4 cbl in2 net29 vdd p12ll_mis_ckt MR=1 L=60n W=120n
XM5 net29 in1 net28 vdd p12ll_mis_ckt MR=1 L=60n W=120n
XM0 net29 qn vss vss n25ll_mis_ckt MR=1 L=280n W=210n
XNM1 vdd q net28 vss n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    cell_PIM2
* View Name:    schematic
************************************************************************

.SUBCKT cell_PIM2 bl cbl in1 in2 sl vdd vss wl
*.PININFO bl:I in1:I in2:I sl:I wl:I cbl:B vdd:B vss:B
XI0 bl q qn sl vdd vss wl / cell_SRAM
XM5 net9 qn vss vss n25ll_mis_ckt MR=1 L=280n W=210n
XM0 net07 qn vss vss n25ll_mis_ckt MR=1 L=280n W=210n
XM3 cbl in2 net9 vdd p12ll_mis_ckt MR=1 L=60n W=120n
XM2 cbl in2 net07 vdd p12ll_mis_ckt MR=1 L=60n W=120n
XM4 net9 in1 net13 vdd p12ll_mis_ckt MR=1 L=60n W=120n
XM1 net07 in1 net7 vdd p12ll_mis_ckt MR=1 L=60n W=120n
XNM3 vdd q net7 vss n12ll_mis_ckt MR=1 L=60n W=120n
XNM4 vdd q net13 vss n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    nand
* View Name:    schematic
************************************************************************

.SUBCKT nand IN0 IN1 OUT VDD VSS
*.PININFO IN0:B IN1:B OUT:B VDD:B VSS:B
XNM4 net10 IN1 VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM3 OUT IN0 net10 VSS n12ll_mis_ckt MR=1 L=60n W=120n
XPM2 OUT IN1 VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM1 OUT IN0 VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv1
* View Name:    schematic
************************************************************************

.SUBCKT inv1 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=60n W=900n
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=60n W=450n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    Tgate
* View Name:    schematic
************************************************************************

.SUBCKT Tgate IN OE OEN OUT VDD VSS
*.PININFO IN:B OE:B OEN:B OUT:B VDD:B VSS:B
XNM2 OUT OE IN VSS n12ll_mis_ckt MR=1 L=60n W=600n
XPM0 IN OEN OUT VDD p12ll_mis_ckt MR=1 L=60n W=1.2u
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    array_test_16r_cell
* View Name:    schematic
************************************************************************

.SUBCKT array_test_16r_cell bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en 
+ in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> in1<9> 
+ in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in2<0> in2<1> in2<2> in2<3> 
+ in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> 
+ in2<14> in2<15> sel sl<0> sl<1> sl<2> sl<3> vdd vss wl<0> wl<1> wl<2> wl<3> 
+ wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15>
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I col_en:I in1<0>:I in1<1>:I in1<2>:I 
*.PININFO in1<3>:I in1<4>:I in1<5>:I in1<6>:I in1<7>:I in1<8>:I in1<9>:I 
*.PININFO in1<10>:I in1<11>:I in1<12>:I in1<13>:I in1<14>:I in1<15>:I in2<0>:I 
*.PININFO in2<1>:I in2<2>:I in2<3>:I in2<4>:I in2<5>:I in2<6>:I in2<7>:I 
*.PININFO in2<8>:I in2<9>:I in2<10>:I in2<11>:I in2<12>:I in2<13>:I in2<14>:I 
*.PININFO in2<15>:I sel:I sl<0>:I sl<1>:I sl<2>:I sl<3>:I wl<0>:I wl<1>:I 
*.PININFO wl<2>:I wl<3>:I wl<4>:I wl<5>:I wl<6>:I wl<7>:I wl<8>:I wl<9>:I 
*.PININFO wl<10>:I wl<11>:I wl<12>:I wl<13>:I wl<14>:I wl<15>:I cbl<0>:B 
*.PININFO cbl<1>:B vdd:B vss:B
XI24707 bl<2> net012 in1<11> in2<11> sl<2> vdd vss wl<11> / cell_PIM
XI24708 bl<2> net012 in1<9> in2<9> sl<2> vdd vss wl<9> / cell_PIM
XI24705 bl<2> net012 in1<10> in2<10> sl<2> vdd vss wl<10> / cell_PIM
XI24709 bl<2> net012 in1<8> in2<8> sl<2> vdd vss wl<8> / cell_PIM
XI24967 bl<2> net012 in1<0> in2<0> sl<2> vdd vss wl<0> / cell_PIM
XI24966 bl<2> net012 in1<1> in2<1> sl<2> vdd vss wl<1> / cell_PIM
XI24965 bl<2> net012 in1<2> in2<2> sl<2> vdd vss wl<2> / cell_PIM
XI24869 bl<2> net012 in1<3> in2<3> sl<2> vdd vss wl<3> / cell_PIM
XI24868 bl<2> net012 in1<4> in2<4> sl<2> vdd vss wl<4> / cell_PIM
XI24867 bl<2> net012 in1<6> in2<6> sl<2> vdd vss wl<6> / cell_PIM
XI24866 bl<2> net012 in1<7> in2<7> sl<2> vdd vss wl<7> / cell_PIM
XI24865 bl<2> net012 in1<5> in2<5> sl<2> vdd vss wl<5> / cell_PIM
XI24698 bl<0> net0145 in1<8> in2<8> sl<0> vdd vss wl<8> / cell_PIM
XI24699 bl<0> net0145 in1<9> in2<9> sl<0> vdd vss wl<9> / cell_PIM
XI24696 bl<0> net0145 in1<11> in2<11> sl<0> vdd vss wl<11> / cell_PIM
XI24695 bl<0> net0145 in1<10> in2<10> sl<0> vdd vss wl<10> / cell_PIM
XI24961 bl<0> net0145 in1<0> in2<0> sl<0> vdd vss wl<0> / cell_PIM
XI24960 bl<0> net0145 in1<2> in2<2> sl<0> vdd vss wl<2> / cell_PIM
XI24959 bl<0> net0145 in1<1> in2<1> sl<0> vdd vss wl<1> / cell_PIM
XI24859 bl<0> net0145 in1<4> in2<4> sl<0> vdd vss wl<4> / cell_PIM
XI24857 bl<0> net0145 in1<7> in2<7> sl<0> vdd vss wl<7> / cell_PIM
XI24856 bl<0> net0145 in1<6> in2<6> sl<0> vdd vss wl<6> / cell_PIM
XI24855 bl<0> net0145 in1<5> in2<5> sl<0> vdd vss wl<5> / cell_PIM
XI24858 bl<0> net0145 in1<3> in2<3> sl<0> vdd vss wl<3> / cell_PIM
XI24706 bl<2> net012 in1<12> in2<12> sl<2> vdd vss wl<12> / cell_PIM
XI24548 bl<2> net012 in1<14> in2<14> sl<2> vdd vss wl<14> / cell_PIM
XI24549 bl<2> net012 in1<13> in2<13> sl<2> vdd vss wl<13> / cell_PIM
XI24545 bl<2> net012 in1<15> in2<15> sl<2> vdd vss wl<15> / cell_PIM
XI24538 bl<0> net0145 in1<13> in2<13> sl<0> vdd vss wl<13> / cell_PIM
XI24697 bl<0> net0145 in1<12> in2<12> sl<0> vdd vss wl<12> / cell_PIM
XI24539 bl<0> net0145 in1<14> in2<14> sl<0> vdd vss wl<14> / cell_PIM
XI24535 bl<0> net0145 in1<15> in2<15> sl<0> vdd vss wl<15> / cell_PIM
XI24711 bl<3> net012 in1<11> in2<11> sl<3> vdd vss wl<11> / cell_PIM2
XI24712 bl<3> net012 in1<10> in2<10> sl<3> vdd vss wl<10> / cell_PIM2
XI24713 bl<3> net012 in1<9> in2<9> sl<3> vdd vss wl<9> / cell_PIM2
XI24970 bl<3> net012 in1<0> in2<0> sl<3> vdd vss wl<0> / cell_PIM2
XI24969 bl<3> net012 in1<1> in2<1> sl<3> vdd vss wl<1> / cell_PIM2
XI24968 bl<3> net012 in1<2> in2<2> sl<3> vdd vss wl<2> / cell_PIM2
XI24874 bl<3> net012 in1<4> in2<4> sl<3> vdd vss wl<4> / cell_PIM2
XI24872 bl<3> net012 in1<5> in2<5> sl<3> vdd vss wl<5> / cell_PIM2
XI24871 bl<3> net012 in1<6> in2<6> sl<3> vdd vss wl<6> / cell_PIM2
XI24870 bl<3> net012 in1<7> in2<7> sl<3> vdd vss wl<7> / cell_PIM2
XI24873 bl<3> net012 in1<3> in2<3> sl<3> vdd vss wl<3> / cell_PIM2
XI24714 bl<3> net012 in1<8> in2<8> sl<3> vdd vss wl<8> / cell_PIM2
XI24704 bl<1> net0145 in1<9> in2<9> sl<1> vdd vss wl<9> / cell_PIM2
XI24703 bl<1> net0145 in1<8> in2<8> sl<1> vdd vss wl<8> / cell_PIM2
XI24701 bl<1> net0145 in1<11> in2<11> sl<1> vdd vss wl<11> / cell_PIM2
XI24700 bl<1> net0145 in1<10> in2<10> sl<1> vdd vss wl<10> / cell_PIM2
XI24964 bl<1> net0145 in1<0> in2<0> sl<1> vdd vss wl<0> / cell_PIM2
XI24962 bl<1> net0145 in1<1> in2<1> sl<1> vdd vss wl<1> / cell_PIM2
XI24963 bl<1> net0145 in1<2> in2<2> sl<1> vdd vss wl<2> / cell_PIM2
XI24864 bl<1> net0145 in1<3> in2<3> sl<1> vdd vss wl<3> / cell_PIM2
XI24862 bl<1> net0145 in1<7> in2<7> sl<1> vdd vss wl<7> / cell_PIM2
XI24861 bl<1> net0145 in1<6> in2<6> sl<1> vdd vss wl<6> / cell_PIM2
XI24860 bl<1> net0145 in1<5> in2<5> sl<1> vdd vss wl<5> / cell_PIM2
XI24863 bl<1> net0145 in1<4> in2<4> sl<1> vdd vss wl<4> / cell_PIM2
XI24710 bl<3> net012 in1<12> in2<12> sl<3> vdd vss wl<12> / cell_PIM2
XI24553 bl<3> net012 in1<14> in2<14> sl<3> vdd vss wl<14> / cell_PIM2
XI24554 bl<3> net012 in1<13> in2<13> sl<3> vdd vss wl<13> / cell_PIM2
XI24552 bl<3> net012 in1<15> in2<15> sl<3> vdd vss wl<15> / cell_PIM2
XI24543 bl<1> net0145 in1<13> in2<13> sl<1> vdd vss wl<13> / cell_PIM2
XI24702 bl<1> net0145 in1<12> in2<12> sl<1> vdd vss wl<12> / cell_PIM2
XI24544 bl<1> net0145 in1<14> in2<14> sl<1> vdd vss wl<14> / cell_PIM2
XI24540 bl<1> net0145 in1<15> in2<15> sl<1> vdd vss wl<15> / cell_PIM2
XI32 sel_n col_en en vdd vss / nand
XI14<0> sel sel_n vdd vss / inv1
XI14<1> sel sel_n vdd vss / inv1
XI14<2> sel sel_n vdd vss / inv1
XI14<3> sel sel_n vdd vss / inv1
XI14<4> sel sel_n vdd vss / inv1
XI14<5> sel sel_n vdd vss / inv1
XI14<6> sel sel_n vdd vss / inv1
XI14<7> sel sel_n vdd vss / inv1
XI14<8> sel sel_n vdd vss / inv1
XI14<9> sel sel_n vdd vss / inv1
XI14<10> sel sel_n vdd vss / inv1
XI14<11> sel sel_n vdd vss / inv1
XI14<12> sel sel_n vdd vss / inv1
XI14<13> sel sel_n vdd vss / inv1
XI14<14> sel sel_n vdd vss / inv1
XI14<15> sel sel_n vdd vss / inv1
XI33<0> en en_n vdd vss / inv1
XI33<1> en en_n vdd vss / inv1
XI33<2> en en_n vdd vss / inv1
XI33<3> en en_n vdd vss / inv1
XI33<4> en en_n vdd vss / inv1
XI33<5> en en_n vdd vss / inv1
XI33<6> en en_n vdd vss / inv1
XI33<7> en en_n vdd vss / inv1
XI33<8> en en_n vdd vss / inv1
XI33<9> en en_n vdd vss / inv1
XI33<10> en en_n vdd vss / inv1
XI33<11> en en_n vdd vss / inv1
XI33<12> en en_n vdd vss / inv1
XI33<13> en en_n vdd vss / inv1
XI33<14> en en_n vdd vss / inv1
XI33<15> en en_n vdd vss / inv1
XI31 net012 en en_n cbl<1> vdd vss / Tgate
XI30 net0145 en en_n cbl<0> vdd vss / Tgate
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    3nand
* View Name:    schematic
************************************************************************

.SUBCKT 3nand VDD VSS in<0> in<1> in<2> out
*.PININFO in<0>:I in<1>:I in<2>:I out:O VDD:B VSS:B
XPM0 out in<0> VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XPM1 out in<2> VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XPM2 out in<1> VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XNM6 net12 in<2> VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
XNM5 net19 in<1> net12 VSS n12ll_mis_ckt MR=1 L=80n W=200n
XNM4 out in<0> net19 VSS n12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv4
* View Name:    schematic
************************************************************************

.SUBCKT inv4 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=60n W=1.8u
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=60n W=3.6u
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    2x4decoder
* View Name:    schematic
************************************************************************

.SUBCKT 2x4decoder VDD VSS en in<0> in<1> nout<0> nout<1> nout<2> nout<3>
*.PININFO en:I in<0>:I in<1>:I nout<0>:O nout<1>:O nout<2>:O nout<3>:O VDD:B 
*.PININFO VSS:B
XI3 VDD VSS in<0> net06 in<1> net016 / 3nand
XI2 VDD VSS net11 net06 in<1> net017 / 3nand
XI1 VDD VSS in<0> net06 net04 net018 / 3nand
XI0 VDD VSS net11 net06 net04 net019 / 3nand
XI6 en net06 VDD VSS / inv1
XI5 in<1> net04 VDD VSS / inv1
XI4 in<0> net11 VDD VSS / inv1
XI44 net016 nout<3> VDD VSS / inv4
XI43 net017 nout<2> VDD VSS / inv4
XI42 net018 nout<1> VDD VSS / inv4
XI41 net019 nout<0> VDD VSS / inv4
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    3x8decoder_2
* View Name:    schematic
************************************************************************

.SUBCKT 3x8decoder_2 en in<0> in<1> in<2> out<0> out<1> out<2> out<3> out<4> 
+ out<5> out<6> out<7> vdd vss
*.PININFO en:I in<0>:I in<1>:I in<2>:I out<0>:O out<1>:O out<2>:O out<3>:O 
*.PININFO out<4>:O out<5>:O out<6>:O out<7>:O vdd:B vss:B
XI1 vdd vss en2 in<0> in<1> out<4> out<5> out<6> out<7> / 2x4decoder
XI0 vdd vss en1 in<0> in<1> out<0> out<1> out<2> out<3> / 2x4decoder
XI6 in<2> en net010 vdd vss / nand
XI7 inn<2> en net09 vdd vss / nand
XI8 net09 en2 vdd vss / inv1
XI5 net010 en1 vdd vss / inv1
XI2 in<2> inn<2> vdd vss / inv1
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    array_test_cel_2
* View Name:    schematic
************************************************************************

.SUBCKT array_test_cel_2 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<0> 
+ in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> 
+ in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> in1<17> in1<18> in1<19> 
+ in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> in1<26> in1<27> in1<28> 
+ in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> in1<35> in1<36> in1<37> 
+ in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> in1<44> in1<45> in1<46> 
+ in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> in1<53> in1<54> in1<55> 
+ in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> in1<62> in1<63> in1<64> 
+ in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> in1<71> in1<72> in1<73> 
+ in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> in1<80> in1<81> in1<82> 
+ in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> in1<89> in1<90> in1<91> 
+ in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> in1<98> in1<99> in1<100> 
+ in1<101> in1<102> in1<103> in1<104> in1<105> in1<106> in1<107> in1<108> 
+ in1<109> in1<110> in1<111> in1<112> in1<113> in1<114> in1<115> in1<116> 
+ in1<117> in1<118> in1<119> in1<120> in1<121> in1<122> in1<123> in1<124> 
+ in1<125> in1<126> in1<127> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> 
+ in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> 
+ in2<17> in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> 
+ in2<26> in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> 
+ in2<35> in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> 
+ in2<44> in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> 
+ in2<53> in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> 
+ in2<62> in2<63> in2<64> in2<65> in2<66> in2<67> in2<68> in2<69> in2<70> 
+ in2<71> in2<72> in2<73> in2<74> in2<75> in2<76> in2<77> in2<78> in2<79> 
+ in2<80> in2<81> in2<82> in2<83> in2<84> in2<85> in2<86> in2<87> in2<88> 
+ in2<89> in2<90> in2<91> in2<92> in2<93> in2<94> in2<95> in2<96> in2<97> 
+ in2<98> in2<99> in2<100> in2<101> in2<102> in2<103> in2<104> in2<105> 
+ in2<106> in2<107> in2<108> in2<109> in2<110> in2<111> in2<112> in2<113> 
+ in2<114> in2<115> in2<116> in2<117> in2<118> in2<119> in2<120> in2<121> 
+ in2<122> in2<123> in2<124> in2<125> in2<126> in2<127> reg_en sel_en sl<0> 
+ sl<1> sl<2> sl<3> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> 
+ wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> 
+ wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> 
+ wl<30> wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> 
+ wl<41> wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> 
+ wl<52> wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> 
+ wl<63> wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> 
+ wl<74> wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> 
+ wl<85> wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> 
+ wl<96> wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> 
+ wl<106> wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> 
+ wl<115> wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> 
+ wl<124> wl<125> wl<126> wl<127>
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I col_en:I in1<0>:I in1<1>:I in1<2>:I 
*.PININFO in1<3>:I in1<4>:I in1<5>:I in1<6>:I in1<7>:I in1<8>:I in1<9>:I 
*.PININFO in1<10>:I in1<11>:I in1<12>:I in1<13>:I in1<14>:I in1<15>:I 
*.PININFO in1<16>:I in1<17>:I in1<18>:I in1<19>:I in1<20>:I in1<21>:I 
*.PININFO in1<22>:I in1<23>:I in1<24>:I in1<25>:I in1<26>:I in1<27>:I 
*.PININFO in1<28>:I in1<29>:I in1<30>:I in1<31>:I in1<32>:I in1<33>:I 
*.PININFO in1<34>:I in1<35>:I in1<36>:I in1<37>:I in1<38>:I in1<39>:I 
*.PININFO in1<40>:I in1<41>:I in1<42>:I in1<43>:I in1<44>:I in1<45>:I 
*.PININFO in1<46>:I in1<47>:I in1<48>:I in1<49>:I in1<50>:I in1<51>:I 
*.PININFO in1<52>:I in1<53>:I in1<54>:I in1<55>:I in1<56>:I in1<57>:I 
*.PININFO in1<58>:I in1<59>:I in1<60>:I in1<61>:I in1<62>:I in1<63>:I 
*.PININFO in1<64>:I in1<65>:I in1<66>:I in1<67>:I in1<68>:I in1<69>:I 
*.PININFO in1<70>:I in1<71>:I in1<72>:I in1<73>:I in1<74>:I in1<75>:I 
*.PININFO in1<76>:I in1<77>:I in1<78>:I in1<79>:I in1<80>:I in1<81>:I 
*.PININFO in1<82>:I in1<83>:I in1<84>:I in1<85>:I in1<86>:I in1<87>:I 
*.PININFO in1<88>:I in1<89>:I in1<90>:I in1<91>:I in1<92>:I in1<93>:I 
*.PININFO in1<94>:I in1<95>:I in1<96>:I in1<97>:I in1<98>:I in1<99>:I 
*.PININFO in1<100>:I in1<101>:I in1<102>:I in1<103>:I in1<104>:I in1<105>:I 
*.PININFO in1<106>:I in1<107>:I in1<108>:I in1<109>:I in1<110>:I in1<111>:I 
*.PININFO in1<112>:I in1<113>:I in1<114>:I in1<115>:I in1<116>:I in1<117>:I 
*.PININFO in1<118>:I in1<119>:I in1<120>:I in1<121>:I in1<122>:I in1<123>:I 
*.PININFO in1<124>:I in1<125>:I in1<126>:I in1<127>:I in2<0>:I in2<1>:I 
*.PININFO in2<2>:I in2<3>:I in2<4>:I in2<5>:I in2<6>:I in2<7>:I in2<8>:I 
*.PININFO in2<9>:I in2<10>:I in2<11>:I in2<12>:I in2<13>:I in2<14>:I in2<15>:I 
*.PININFO in2<16>:I in2<17>:I in2<18>:I in2<19>:I in2<20>:I in2<21>:I 
*.PININFO in2<22>:I in2<23>:I in2<24>:I in2<25>:I in2<26>:I in2<27>:I 
*.PININFO in2<28>:I in2<29>:I in2<30>:I in2<31>:I in2<32>:I in2<33>:I 
*.PININFO in2<34>:I in2<35>:I in2<36>:I in2<37>:I in2<38>:I in2<39>:I 
*.PININFO in2<40>:I in2<41>:I in2<42>:I in2<43>:I in2<44>:I in2<45>:I 
*.PININFO in2<46>:I in2<47>:I in2<48>:I in2<49>:I in2<50>:I in2<51>:I 
*.PININFO in2<52>:I in2<53>:I in2<54>:I in2<55>:I in2<56>:I in2<57>:I 
*.PININFO in2<58>:I in2<59>:I in2<60>:I in2<61>:I in2<62>:I in2<63>:I 
*.PININFO in2<64>:I in2<65>:I in2<66>:I in2<67>:I in2<68>:I in2<69>:I 
*.PININFO in2<70>:I in2<71>:I in2<72>:I in2<73>:I in2<74>:I in2<75>:I 
*.PININFO in2<76>:I in2<77>:I in2<78>:I in2<79>:I in2<80>:I in2<81>:I 
*.PININFO in2<82>:I in2<83>:I in2<84>:I in2<85>:I in2<86>:I in2<87>:I 
*.PININFO in2<88>:I in2<89>:I in2<90>:I in2<91>:I in2<92>:I in2<93>:I 
*.PININFO in2<94>:I in2<95>:I in2<96>:I in2<97>:I in2<98>:I in2<99>:I 
*.PININFO in2<100>:I in2<101>:I in2<102>:I in2<103>:I in2<104>:I in2<105>:I 
*.PININFO in2<106>:I in2<107>:I in2<108>:I in2<109>:I in2<110>:I in2<111>:I 
*.PININFO in2<112>:I in2<113>:I in2<114>:I in2<115>:I in2<116>:I in2<117>:I 
*.PININFO in2<118>:I in2<119>:I in2<120>:I in2<121>:I in2<122>:I in2<123>:I 
*.PININFO in2<124>:I in2<125>:I in2<126>:I in2<127>:I reg_en:I sel_en:I 
*.PININFO sl<0>:I sl<1>:I sl<2>:I sl<3>:I wl<0>:I wl<1>:I wl<2>:I wl<3>:I 
*.PININFO wl<4>:I wl<5>:I wl<6>:I wl<7>:I wl<8>:I wl<9>:I wl<10>:I wl<11>:I 
*.PININFO wl<12>:I wl<13>:I wl<14>:I wl<15>:I wl<16>:I wl<17>:I wl<18>:I 
*.PININFO wl<19>:I wl<20>:I wl<21>:I wl<22>:I wl<23>:I wl<24>:I wl<25>:I 
*.PININFO wl<26>:I wl<27>:I wl<28>:I wl<29>:I wl<30>:I wl<31>:I wl<32>:I 
*.PININFO wl<33>:I wl<34>:I wl<35>:I wl<36>:I wl<37>:I wl<38>:I wl<39>:I 
*.PININFO wl<40>:I wl<41>:I wl<42>:I wl<43>:I wl<44>:I wl<45>:I wl<46>:I 
*.PININFO wl<47>:I wl<48>:I wl<49>:I wl<50>:I wl<51>:I wl<52>:I wl<53>:I 
*.PININFO wl<54>:I wl<55>:I wl<56>:I wl<57>:I wl<58>:I wl<59>:I wl<60>:I 
*.PININFO wl<61>:I wl<62>:I wl<63>:I wl<64>:I wl<65>:I wl<66>:I wl<67>:I 
*.PININFO wl<68>:I wl<69>:I wl<70>:I wl<71>:I wl<72>:I wl<73>:I wl<74>:I 
*.PININFO wl<75>:I wl<76>:I wl<77>:I wl<78>:I wl<79>:I wl<80>:I wl<81>:I 
*.PININFO wl<82>:I wl<83>:I wl<84>:I wl<85>:I wl<86>:I wl<87>:I wl<88>:I 
*.PININFO wl<89>:I wl<90>:I wl<91>:I wl<92>:I wl<93>:I wl<94>:I wl<95>:I 
*.PININFO wl<96>:I wl<97>:I wl<98>:I wl<99>:I wl<100>:I wl<101>:I wl<102>:I 
*.PININFO wl<103>:I wl<104>:I wl<105>:I wl<106>:I wl<107>:I wl<108>:I 
*.PININFO wl<109>:I wl<110>:I wl<111>:I wl<112>:I wl<113>:I wl<114>:I 
*.PININFO wl<115>:I wl<116>:I wl<117>:I wl<118>:I wl<119>:I wl<120>:I 
*.PININFO wl<121>:I wl<122>:I wl<123>:I wl<124>:I wl<125>:I wl<126>:I 
*.PININFO wl<127>:I cbl<0>:O cbl<1>:O vdd:B vss:B
XI25097 bl<2> cbl<1> vdd vdd sl<2> vdd vss vss / cell_PIM
XI25095 bl<0> cbl<0> vdd vdd sl<0> vdd vss vss / cell_PIM
XI49 bl<0> cbl<0> vdd vdd sl<0> vdd vss vss / cell_PIM
XI36 bl<2> cbl<1> vdd vdd sl<2> vdd vss vss / cell_PIM
XI25098 bl<3> cbl<1> vdd vdd sl<3> vdd vss vss / cell_PIM2
XI83 bl<1> cbl<0> vdd vdd sl<1> vdd vss vss / cell_PIM2
XI25096 bl<1> cbl<0> vdd vdd sl<1> vdd vss vss / cell_PIM2
XI69 bl<3> cbl<1> vdd vdd sl<3> vdd vss vss / cell_PIM2
XI117 reg_en sel_en net021 vdd vss / nand
XI114 bl<2> net058 q<2> sl<2> vdd vss wl_reg / cell_SRAM
XI113 bl<1> net059 q<1> sl<1> vdd vss wl_reg / cell_SRAM
XI0 bl<0> net060 q<0> sl<0> vdd vss wl_reg / cell_SRAM
XI112 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<112> in1<113> in1<114> 
+ in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> in1<122> 
+ in1<123> in1<124> in1<125> in1<126> in1<127> in2<112> in2<113> in2<114> 
+ in2<115> in2<116> in2<117> in2<118> in2<119> in2<120> in2<121> in2<122> 
+ in2<123> in2<124> in2<125> in2<126> in2<127> sel<7> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<112> wl<113> wl<114> wl<115> wl<116> wl<117> wl<118> wl<119> 
+ wl<120> wl<121> wl<122> wl<123> wl<124> wl<125> wl<126> wl<127> / 
+ array_test_16r_cell
XI111 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<96> in1<97> in1<98> 
+ in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> in1<106> 
+ in1<107> in1<108> in1<109> in1<110> in1<111> in2<96> in2<97> in2<98> in2<99> 
+ in2<100> in2<101> in2<102> in2<103> in2<104> in2<105> in2<106> in2<107> 
+ in2<108> in2<109> in2<110> in2<111> sel<6> sl<0> sl<1> sl<2> sl<3> vdd vss 
+ wl<96> wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> 
+ wl<106> wl<107> wl<108> wl<109> wl<110> wl<111> / array_test_16r_cell
XI110 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<80> in1<81> in1<82> 
+ in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> in1<89> in1<90> in1<91> 
+ in1<92> in1<93> in1<94> in1<95> in2<80> in2<81> in2<82> in2<83> in2<84> 
+ in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> 
+ in2<94> in2<95> sel<5> sl<0> sl<1> sl<2> sl<3> vdd vss wl<80> wl<81> wl<82> 
+ wl<83> wl<84> wl<85> wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> 
+ wl<94> wl<95> / array_test_16r_cell
XI109 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<64> in1<65> in1<66> 
+ in1<67> in1<68> in1<69> in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> 
+ in1<76> in1<77> in1<78> in1<79> in2<64> in2<65> in2<66> in2<67> in2<68> 
+ in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> in2<76> in2<77> 
+ in2<78> in2<79> sel<4> sl<0> sl<1> sl<2> sl<3> vdd vss wl<64> wl<65> wl<66> 
+ wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> wl<75> wl<76> wl<77> 
+ wl<78> wl<79> / array_test_16r_cell
XI108 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<48> in1<49> in1<50> 
+ in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> 
+ in1<60> in1<61> in1<62> in1<63> in2<48> in2<49> in2<50> in2<51> in2<52> 
+ in2<53> in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> 
+ in2<62> in2<63> sel<3> sl<0> sl<1> sl<2> sl<3> vdd vss wl<48> wl<49> wl<50> 
+ wl<51> wl<52> wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> 
+ wl<62> wl<63> / array_test_16r_cell
XI107 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<32> in1<33> in1<34> 
+ in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> 
+ in1<44> in1<45> in1<46> in1<47> in2<32> in2<33> in2<34> in2<35> in2<36> 
+ in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> 
+ in2<46> in2<47> sel<2> sl<0> sl<1> sl<2> sl<3> vdd vss wl<32> wl<33> wl<34> 
+ wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> wl<42> wl<43> wl<44> wl<45> 
+ wl<46> wl<47> / array_test_16r_cell
XI106 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<16> in1<17> in1<18> 
+ in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> in1<26> in1<27> 
+ in1<28> in1<29> in1<30> in1<31> in2<16> in2<17> in2<18> in2<19> in2<20> 
+ in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> 
+ in2<30> in2<31> sel<1> sl<0> sl<1> sl<2> sl<3> vdd vss wl<16> wl<17> wl<18> 
+ wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> 
+ wl<30> wl<31> / array_test_16r_cell
XI105 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<0> in1<1> in1<2> in1<3> 
+ in1<4> in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> 
+ in1<14> in1<15> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> 
+ in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> sel<0> sl<0> 
+ sl<1> sl<2> sl<3> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> 
+ wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> / array_test_16r_cell
XI116 col_en q<0> q<1> q<2> sel<0> sel<1> sel<2> sel<3> sel<4> sel<5> sel<6> 
+ sel<7> vdd vss / 3x8decoder_2
XI118 net021 wl_reg vdd vss / inv1
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    array_test
* View Name:    schematic
************************************************************************

.SUBCKT array_test bl<0> bl<1> bl<2> bl<3> bl<4> bl<5> bl<6> bl<7> bl<8> bl<9> 
+ bl<10> bl<11> bl<12> bl<13> bl<14> bl<15> bl<16> bl<17> bl<18> bl<19> bl<20> 
+ bl<21> bl<22> bl<23> bl<24> bl<25> bl<26> bl<27> bl<28> bl<29> bl<30> bl<31> 
+ bl<32> bl<33> bl<34> bl<35> bl<36> bl<37> bl<38> bl<39> bl<40> bl<41> bl<42> 
+ bl<43> bl<44> bl<45> bl<46> bl<47> bl<48> bl<49> bl<50> bl<51> bl<52> bl<53> 
+ bl<54> bl<55> bl<56> bl<57> bl<58> bl<59> bl<60> bl<61> bl<62> bl<63> cbl<0> 
+ cbl<1> cbl<2> cbl<3> cbl<4> cbl<5> cbl<6> cbl<7> cbl<8> cbl<9> cbl<10> 
+ cbl<11> cbl<12> cbl<13> cbl<14> cbl<15> cbl<16> cbl<17> cbl<18> cbl<19> 
+ cbl<20> cbl<21> cbl<22> cbl<23> cbl<24> cbl<25> cbl<26> cbl<27> cbl<28> 
+ cbl<29> cbl<30> cbl<31> col_en in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> 
+ in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> 
+ in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> 
+ in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> 
+ in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> 
+ in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> 
+ in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> 
+ in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> 
+ in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> 
+ in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> 
+ in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> 
+ in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> 
+ in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> 
+ in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> 
+ in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> 
+ in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> 
+ in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> 
+ in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> 
+ in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> 
+ in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> 
+ in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> 
+ in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> 
+ in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> 
+ in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> 
+ in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> 
+ in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> 
+ in2<102> in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> 
+ in2<110> in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> 
+ in2<118> in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> 
+ in2<126> in2<127> reg_en sel<0> sel<1> sel<2> sel<3> sel<4> sel<5> sel<6> 
+ sel<7> sel<8> sel<9> sel<10> sel<11> sel<12> sel<13> sel<14> sel<15> sl<0> 
+ sl<1> sl<2> sl<3> sl<4> sl<5> sl<6> sl<7> sl<8> sl<9> sl<10> sl<11> sl<12> 
+ sl<13> sl<14> sl<15> sl<16> sl<17> sl<18> sl<19> sl<20> sl<21> sl<22> sl<23> 
+ sl<24> sl<25> sl<26> sl<27> sl<28> sl<29> sl<30> sl<31> sl<32> sl<33> sl<34> 
+ sl<35> sl<36> sl<37> sl<38> sl<39> sl<40> sl<41> sl<42> sl<43> sl<44> sl<45> 
+ sl<46> sl<47> sl<48> sl<49> sl<50> sl<51> sl<52> sl<53> sl<54> sl<55> sl<56> 
+ sl<57> sl<58> sl<59> sl<60> sl<61> sl<62> sl<63> vdd vss wl<0> wl<1> wl<2> 
+ wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> 
+ wl<15> wl<16> wl<17> wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> 
+ wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> 
+ wl<37> wl<38> wl<39> wl<40> wl<41> wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> 
+ wl<48> wl<49> wl<50> wl<51> wl<52> wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> 
+ wl<59> wl<60> wl<61> wl<62> wl<63> wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> 
+ wl<70> wl<71> wl<72> wl<73> wl<74> wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> 
+ wl<81> wl<82> wl<83> wl<84> wl<85> wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> 
+ wl<92> wl<93> wl<94> wl<95> wl<96> wl<97> wl<98> wl<99> wl<100> wl<101> 
+ wl<102> wl<103> wl<104> wl<105> wl<106> wl<107> wl<108> wl<109> wl<110> 
+ wl<111> wl<112> wl<113> wl<114> wl<115> wl<116> wl<117> wl<118> wl<119> 
+ wl<120> wl<121> wl<122> wl<123> wl<124> wl<125> wl<126> wl<127>
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I bl<4>:I bl<5>:I bl<6>:I bl<7>:I 
*.PININFO bl<8>:I bl<9>:I bl<10>:I bl<11>:I bl<12>:I bl<13>:I bl<14>:I 
*.PININFO bl<15>:I bl<16>:I bl<17>:I bl<18>:I bl<19>:I bl<20>:I bl<21>:I 
*.PININFO bl<22>:I bl<23>:I bl<24>:I bl<25>:I bl<26>:I bl<27>:I bl<28>:I 
*.PININFO bl<29>:I bl<30>:I bl<31>:I bl<32>:I bl<33>:I bl<34>:I bl<35>:I 
*.PININFO bl<36>:I bl<37>:I bl<38>:I bl<39>:I bl<40>:I bl<41>:I bl<42>:I 
*.PININFO bl<43>:I bl<44>:I bl<45>:I bl<46>:I bl<47>:I bl<48>:I bl<49>:I 
*.PININFO bl<50>:I bl<51>:I bl<52>:I bl<53>:I bl<54>:I bl<55>:I bl<56>:I 
*.PININFO bl<57>:I bl<58>:I bl<59>:I bl<60>:I bl<61>:I bl<62>:I bl<63>:I 
*.PININFO col_en:I in1<0>:I in1<1>:I in1<2>:I in1<3>:I in1<4>:I in1<5>:I 
*.PININFO in1<6>:I in1<7>:I in1<8>:I in1<9>:I in1<10>:I in1<11>:I in1<12>:I 
*.PININFO in1<13>:I in1<14>:I in1<15>:I in1<16>:I in1<17>:I in1<18>:I 
*.PININFO in1<19>:I in1<20>:I in1<21>:I in1<22>:I in1<23>:I in1<24>:I 
*.PININFO in1<25>:I in1<26>:I in1<27>:I in1<28>:I in1<29>:I in1<30>:I 
*.PININFO in1<31>:I in1<32>:I in1<33>:I in1<34>:I in1<35>:I in1<36>:I 
*.PININFO in1<37>:I in1<38>:I in1<39>:I in1<40>:I in1<41>:I in1<42>:I 
*.PININFO in1<43>:I in1<44>:I in1<45>:I in1<46>:I in1<47>:I in1<48>:I 
*.PININFO in1<49>:I in1<50>:I in1<51>:I in1<52>:I in1<53>:I in1<54>:I 
*.PININFO in1<55>:I in1<56>:I in1<57>:I in1<58>:I in1<59>:I in1<60>:I 
*.PININFO in1<61>:I in1<62>:I in1<63>:I in1<64>:I in1<65>:I in1<66>:I 
*.PININFO in1<67>:I in1<68>:I in1<69>:I in1<70>:I in1<71>:I in1<72>:I 
*.PININFO in1<73>:I in1<74>:I in1<75>:I in1<76>:I in1<77>:I in1<78>:I 
*.PININFO in1<79>:I in1<80>:I in1<81>:I in1<82>:I in1<83>:I in1<84>:I 
*.PININFO in1<85>:I in1<86>:I in1<87>:I in1<88>:I in1<89>:I in1<90>:I 
*.PININFO in1<91>:I in1<92>:I in1<93>:I in1<94>:I in1<95>:I in1<96>:I 
*.PININFO in1<97>:I in1<98>:I in1<99>:I in1<100>:I in1<101>:I in1<102>:I 
*.PININFO in1<103>:I in1<104>:I in1<105>:I in1<106>:I in1<107>:I in1<108>:I 
*.PININFO in1<109>:I in1<110>:I in1<111>:I in1<112>:I in1<113>:I in1<114>:I 
*.PININFO in1<115>:I in1<116>:I in1<117>:I in1<118>:I in1<119>:I in1<120>:I 
*.PININFO in1<121>:I in1<122>:I in1<123>:I in1<124>:I in1<125>:I in1<126>:I 
*.PININFO in1<127>:I in2<0>:I in2<1>:I in2<2>:I in2<3>:I in2<4>:I in2<5>:I 
*.PININFO in2<6>:I in2<7>:I in2<8>:I in2<9>:I in2<10>:I in2<11>:I in2<12>:I 
*.PININFO in2<13>:I in2<14>:I in2<15>:I in2<16>:I in2<17>:I in2<18>:I 
*.PININFO in2<19>:I in2<20>:I in2<21>:I in2<22>:I in2<23>:I in2<24>:I 
*.PININFO in2<25>:I in2<26>:I in2<27>:I in2<28>:I in2<29>:I in2<30>:I 
*.PININFO in2<31>:I in2<32>:I in2<33>:I in2<34>:I in2<35>:I in2<36>:I 
*.PININFO in2<37>:I in2<38>:I in2<39>:I in2<40>:I in2<41>:I in2<42>:I 
*.PININFO in2<43>:I in2<44>:I in2<45>:I in2<46>:I in2<47>:I in2<48>:I 
*.PININFO in2<49>:I in2<50>:I in2<51>:I in2<52>:I in2<53>:I in2<54>:I 
*.PININFO in2<55>:I in2<56>:I in2<57>:I in2<58>:I in2<59>:I in2<60>:I 
*.PININFO in2<61>:I in2<62>:I in2<63>:I in2<64>:I in2<65>:I in2<66>:I 
*.PININFO in2<67>:I in2<68>:I in2<69>:I in2<70>:I in2<71>:I in2<72>:I 
*.PININFO in2<73>:I in2<74>:I in2<75>:I in2<76>:I in2<77>:I in2<78>:I 
*.PININFO in2<79>:I in2<80>:I in2<81>:I in2<82>:I in2<83>:I in2<84>:I 
*.PININFO in2<85>:I in2<86>:I in2<87>:I in2<88>:I in2<89>:I in2<90>:I 
*.PININFO in2<91>:I in2<92>:I in2<93>:I in2<94>:I in2<95>:I in2<96>:I 
*.PININFO in2<97>:I in2<98>:I in2<99>:I in2<100>:I in2<101>:I in2<102>:I 
*.PININFO in2<103>:I in2<104>:I in2<105>:I in2<106>:I in2<107>:I in2<108>:I 
*.PININFO in2<109>:I in2<110>:I in2<111>:I in2<112>:I in2<113>:I in2<114>:I 
*.PININFO in2<115>:I in2<116>:I in2<117>:I in2<118>:I in2<119>:I in2<120>:I 
*.PININFO in2<121>:I in2<122>:I in2<123>:I in2<124>:I in2<125>:I in2<126>:I 
*.PININFO in2<127>:I reg_en:I sel<0>:I sel<1>:I sel<2>:I sel<3>:I sel<4>:I 
*.PININFO sel<5>:I sel<6>:I sel<7>:I sel<8>:I sel<9>:I sel<10>:I sel<11>:I 
*.PININFO sel<12>:I sel<13>:I sel<14>:I sel<15>:I sl<0>:I sl<1>:I sl<2>:I 
*.PININFO sl<3>:I sl<4>:I sl<5>:I sl<6>:I sl<7>:I sl<8>:I sl<9>:I sl<10>:I 
*.PININFO sl<11>:I sl<12>:I sl<13>:I sl<14>:I sl<15>:I sl<16>:I sl<17>:I 
*.PININFO sl<18>:I sl<19>:I sl<20>:I sl<21>:I sl<22>:I sl<23>:I sl<24>:I 
*.PININFO sl<25>:I sl<26>:I sl<27>:I sl<28>:I sl<29>:I sl<30>:I sl<31>:I 
*.PININFO sl<32>:I sl<33>:I sl<34>:I sl<35>:I sl<36>:I sl<37>:I sl<38>:I 
*.PININFO sl<39>:I sl<40>:I sl<41>:I sl<42>:I sl<43>:I sl<44>:I sl<45>:I 
*.PININFO sl<46>:I sl<47>:I sl<48>:I sl<49>:I sl<50>:I sl<51>:I sl<52>:I 
*.PININFO sl<53>:I sl<54>:I sl<55>:I sl<56>:I sl<57>:I sl<58>:I sl<59>:I 
*.PININFO sl<60>:I sl<61>:I sl<62>:I sl<63>:I wl<0>:I wl<1>:I wl<2>:I wl<3>:I 
*.PININFO wl<4>:I wl<5>:I wl<6>:I wl<7>:I wl<8>:I wl<9>:I wl<10>:I wl<11>:I 
*.PININFO wl<12>:I wl<13>:I wl<14>:I wl<15>:I wl<16>:I wl<17>:I wl<18>:I 
*.PININFO wl<19>:I wl<20>:I wl<21>:I wl<22>:I wl<23>:I wl<24>:I wl<25>:I 
*.PININFO wl<26>:I wl<27>:I wl<28>:I wl<29>:I wl<30>:I wl<31>:I wl<32>:I 
*.PININFO wl<33>:I wl<34>:I wl<35>:I wl<36>:I wl<37>:I wl<38>:I wl<39>:I 
*.PININFO wl<40>:I wl<41>:I wl<42>:I wl<43>:I wl<44>:I wl<45>:I wl<46>:I 
*.PININFO wl<47>:I wl<48>:I wl<49>:I wl<50>:I wl<51>:I wl<52>:I wl<53>:I 
*.PININFO wl<54>:I wl<55>:I wl<56>:I wl<57>:I wl<58>:I wl<59>:I wl<60>:I 
*.PININFO wl<61>:I wl<62>:I wl<63>:I wl<64>:I wl<65>:I wl<66>:I wl<67>:I 
*.PININFO wl<68>:I wl<69>:I wl<70>:I wl<71>:I wl<72>:I wl<73>:I wl<74>:I 
*.PININFO wl<75>:I wl<76>:I wl<77>:I wl<78>:I wl<79>:I wl<80>:I wl<81>:I 
*.PININFO wl<82>:I wl<83>:I wl<84>:I wl<85>:I wl<86>:I wl<87>:I wl<88>:I 
*.PININFO wl<89>:I wl<90>:I wl<91>:I wl<92>:I wl<93>:I wl<94>:I wl<95>:I 
*.PININFO wl<96>:I wl<97>:I wl<98>:I wl<99>:I wl<100>:I wl<101>:I wl<102>:I 
*.PININFO wl<103>:I wl<104>:I wl<105>:I wl<106>:I wl<107>:I wl<108>:I 
*.PININFO wl<109>:I wl<110>:I wl<111>:I wl<112>:I wl<113>:I wl<114>:I 
*.PININFO wl<115>:I wl<116>:I wl<117>:I wl<118>:I wl<119>:I wl<120>:I 
*.PININFO wl<121>:I wl<122>:I wl<123>:I wl<124>:I wl<125>:I wl<126>:I 
*.PININFO wl<127>:I cbl<0>:O cbl<1>:O cbl<2>:O cbl<3>:O cbl<4>:O cbl<5>:O 
*.PININFO cbl<6>:O cbl<7>:O cbl<8>:O cbl<9>:O cbl<10>:O cbl<11>:O cbl<12>:O 
*.PININFO cbl<13>:O cbl<14>:O cbl<15>:O cbl<16>:O cbl<17>:O cbl<18>:O 
*.PININFO cbl<19>:O cbl<20>:O cbl<21>:O cbl<22>:O cbl<23>:O cbl<24>:O 
*.PININFO cbl<25>:O cbl<26>:O cbl<27>:O cbl<28>:O cbl<29>:O cbl<30>:O 
*.PININFO cbl<31>:O vdd:B vss:B
XI25357 vss vss in1<0> in2<0> vss vdd vss wl<0> / cell_PIM
XI25358 vss vss vdd vdd vss vdd vss vss / cell_PIM
XI25354 vss vss in1<4> in2<4> vss vdd vss wl<4> / cell_PIM
XI25355 vss vss in1<1> in2<1> vss vdd vss wl<1> / cell_PIM
XI25356 vss vss in1<2> in2<2> vss vdd vss wl<2> / cell_PIM
XI25352 vss vss in1<7> in2<7> vss vdd vss wl<7> / cell_PIM
XI25351 vss vss in1<6> in2<6> vss vdd vss wl<6> / cell_PIM
XI25350 vss vss in1<5> in2<5> vss vdd vss wl<5> / cell_PIM
XI25349 vss vss in1<9> in2<9> vss vdd vss wl<9> / cell_PIM
XI25353 vss vss in1<3> in2<3> vss vdd vss wl<3> / cell_PIM
XI25348 vss vss in1<8> in2<8> vss vdd vss wl<8> / cell_PIM
XI25347 vss vss in1<11> in2<11> vss vdd vss wl<11> / cell_PIM
XI25346 vss vss in1<10> in2<10> vss vdd vss wl<10> / cell_PIM
XI25345 vss vss in1<12> in2<12> vss vdd vss wl<12> / cell_PIM
XI25344 vss vss in1<14> in2<14> vss vdd vss wl<14> / cell_PIM
XI25342 vss vss in1<16> in2<16> vss vdd vss wl<16> / cell_PIM
XI25341 vss vss in1<15> in2<15> vss vdd vss wl<15> / cell_PIM
XI25340 vss vss in1<17> in2<17> vss vdd vss wl<17> / cell_PIM
XI25339 vss vss in1<19> in2<19> vss vdd vss wl<19> / cell_PIM
XI25343 vss vss in1<13> in2<13> vss vdd vss wl<13> / cell_PIM
XI25337 vss vss in1<21> in2<21> vss vdd vss wl<21> / cell_PIM
XI25336 vss vss in1<20> in2<20> vss vdd vss wl<20> / cell_PIM
XI25335 vss vss in1<24> in2<24> vss vdd vss wl<24> / cell_PIM
XI25334 vss vss in1<23> in2<23> vss vdd vss wl<23> / cell_PIM
XI25338 vss vss in1<18> in2<18> vss vdd vss wl<18> / cell_PIM
XI25332 vss vss in1<26> in2<26> vss vdd vss wl<26> / cell_PIM
XI25331 vss vss in1<25> in2<25> vss vdd vss wl<25> / cell_PIM
XI25330 vss vss in1<28> in2<28> vss vdd vss wl<28> / cell_PIM
XI25329 vss vss in1<27> in2<27> vss vdd vss wl<27> / cell_PIM
XI25333 vss vss in1<22> in2<22> vss vdd vss wl<22> / cell_PIM
XI25328 vss vss in1<31> in2<31> vss vdd vss wl<31> / cell_PIM
XI25327 vss vss in1<30> in2<30> vss vdd vss wl<30> / cell_PIM
XI25326 vss vss in1<29> in2<29> vss vdd vss wl<29> / cell_PIM
XI25325 vss vss in1<33> in2<33> vss vdd vss wl<33> / cell_PIM
XI25324 vss vss in1<32> in2<32> vss vdd vss wl<32> / cell_PIM
XI25322 vss vss in1<34> in2<34> vss vdd vss wl<34> / cell_PIM
XI25321 vss vss in1<36> in2<36> vss vdd vss wl<36> / cell_PIM
XI25320 vss vss in1<38> in2<38> vss vdd vss wl<38> / cell_PIM
XI25319 vss vss in1<37> in2<37> vss vdd vss wl<37> / cell_PIM
XI25323 vss vss in1<35> in2<35> vss vdd vss wl<35> / cell_PIM
XI25317 vss vss in1<39> in2<39> vss vdd vss wl<39> / cell_PIM
XI25316 vss vss in1<41> in2<41> vss vdd vss wl<41> / cell_PIM
XI25315 vss vss in1<43> in2<43> vss vdd vss wl<43> / cell_PIM
XI25314 vss vss in1<42> in2<42> vss vdd vss wl<42> / cell_PIM
XI25318 vss vss in1<40> in2<40> vss vdd vss wl<40> / cell_PIM
XI25312 vss vss in1<44> in2<44> vss vdd vss wl<44> / cell_PIM
XI25311 vss vss in1<47> in2<47> vss vdd vss wl<47> / cell_PIM
XI25310 vss vss in1<46> in2<46> vss vdd vss wl<46> / cell_PIM
XI25309 vss vss in1<50> in2<50> vss vdd vss wl<50> / cell_PIM
XI25313 vss vss in1<45> in2<45> vss vdd vss wl<45> / cell_PIM
XI25308 vss vss in1<49> in2<49> vss vdd vss wl<49> / cell_PIM
XI25307 vss vss in1<48> in2<48> vss vdd vss wl<48> / cell_PIM
XI25306 vss vss in1<52> in2<52> vss vdd vss wl<52> / cell_PIM
XI25305 vss vss in1<51> in2<51> vss vdd vss wl<51> / cell_PIM
XI25304 vss vss in1<55> in2<55> vss vdd vss wl<55> / cell_PIM
XI25302 vss vss in1<53> in2<53> vss vdd vss wl<53> / cell_PIM
XI25301 vss vss in1<57> in2<57> vss vdd vss wl<57> / cell_PIM
XI25300 vss vss in1<56> in2<56> vss vdd vss wl<56> / cell_PIM
XI25299 vss vss in1<59> in2<59> vss vdd vss wl<59> / cell_PIM
XI25303 vss vss in1<54> in2<54> vss vdd vss wl<54> / cell_PIM
XI25297 vss vss in1<60> in2<60> vss vdd vss wl<60> / cell_PIM
XI25296 vss vss in1<62> in2<62> vss vdd vss wl<62> / cell_PIM
XI25295 vss vss in1<61> in2<61> vss vdd vss wl<61> / cell_PIM
XI25294 vss vss in1<64> in2<64> vss vdd vss wl<64> / cell_PIM
XI25298 vss vss in1<58> in2<58> vss vdd vss wl<58> / cell_PIM
XI25292 vss vss in1<65> in2<65> vss vdd vss wl<65> / cell_PIM
XI25291 vss vss in1<67> in2<67> vss vdd vss wl<67> / cell_PIM
XI25290 vss vss in1<66> in2<66> vss vdd vss wl<66> / cell_PIM
XI25289 vss vss in1<69> in2<69> vss vdd vss wl<69> / cell_PIM
XI25293 vss vss in1<63> in2<63> vss vdd vss wl<63> / cell_PIM
XI25288 vss vss in1<68> in2<68> vss vdd vss wl<68> / cell_PIM
XI25287 vss vss in1<70> in2<70> vss vdd vss wl<70> / cell_PIM
XI25286 vss vss in1<71> in2<71> vss vdd vss wl<71> / cell_PIM
XI25285 vss vss in1<74> in2<74> vss vdd vss wl<74> / cell_PIM
XI25284 vss vss in1<73> in2<73> vss vdd vss wl<73> / cell_PIM
XI25282 vss vss in1<75> in2<75> vss vdd vss wl<75> / cell_PIM
XI25281 vss vss in1<76> in2<76> vss vdd vss wl<76> / cell_PIM
XI25280 vss vss in1<79> in2<79> vss vdd vss wl<79> / cell_PIM
XI25279 vss vss in1<78> in2<78> vss vdd vss wl<78> / cell_PIM
XI25283 vss vss in1<72> in2<72> vss vdd vss wl<72> / cell_PIM
XI25277 vss vss in1<80> in2<80> vss vdd vss wl<80> / cell_PIM
XI25276 vss vss in1<81> in2<81> vss vdd vss wl<81> / cell_PIM
XI25275 vss vss in1<83> in2<83> vss vdd vss wl<83> / cell_PIM
XI25274 vss vss in1<82> in2<82> vss vdd vss wl<82> / cell_PIM
XI25278 vss vss in1<77> in2<77> vss vdd vss wl<77> / cell_PIM
XI25272 vss vss in1<86> in2<86> vss vdd vss wl<86> / cell_PIM
XI25271 vss vss in1<85> in2<85> vss vdd vss wl<85> / cell_PIM
XI25270 vss vss in1<88> in2<88> vss vdd vss wl<88> / cell_PIM
XI25269 vss vss in1<87> in2<87> vss vdd vss wl<87> / cell_PIM
XI25273 vss vss in1<84> in2<84> vss vdd vss wl<84> / cell_PIM
XI25268 vss vss in1<89> in2<89> vss vdd vss wl<89> / cell_PIM
XI25267 vss vss in1<91> in2<91> vss vdd vss wl<91> / cell_PIM
XI25266 vss vss in1<90> in2<90> vss vdd vss wl<90> / cell_PIM
XI25265 vss vss in1<93> in2<93> vss vdd vss wl<93> / cell_PIM
XI25264 vss vss in1<92> in2<92> vss vdd vss wl<92> / cell_PIM
XI25262 vss vss in1<95> in2<95> vss vdd vss wl<95> / cell_PIM
XI25261 vss vss in1<98> in2<98> vss vdd vss wl<98> / cell_PIM
XI25260 vss vss in1<97> in2<97> vss vdd vss wl<97> / cell_PIM
XI25259 vss vss in1<96> in2<96> vss vdd vss wl<96> / cell_PIM
XI25263 vss vss in1<94> in2<94> vss vdd vss wl<94> / cell_PIM
XI25257 vss vss in1<100> in2<100> vss vdd vss wl<100> / cell_PIM
XI25256 vss vss in1<103> in2<103> vss vdd vss wl<103> / cell_PIM
XI25255 vss vss in1<102> in2<102> vss vdd vss wl<102> / cell_PIM
XI25254 vss vss in1<101> in2<101> vss vdd vss wl<101> / cell_PIM
XI25258 vss vss in1<99> in2<99> vss vdd vss wl<99> / cell_PIM
XI25252 vss vss in1<105> in2<105> vss vdd vss wl<105> / cell_PIM
XI25251 vss vss in1<107> in2<107> vss vdd vss wl<107> / cell_PIM
XI25250 vss vss in1<106> in2<106> vss vdd vss wl<106> / cell_PIM
XI25249 vss vss in1<108> in2<108> vss vdd vss wl<108> / cell_PIM
XI25253 vss vss in1<104> in2<104> vss vdd vss wl<104> / cell_PIM
XI25248 vss vss in1<109> in2<109> vss vdd vss wl<109> / cell_PIM
XI25247 vss vss in1<110> in2<110> vss vdd vss wl<110> / cell_PIM
XI25246 vss vss in1<112> in2<112> vss vdd vss wl<112> / cell_PIM
XI25245 vss vss in1<111> in2<111> vss vdd vss wl<111> / cell_PIM
XI25244 vss vss in1<113> in2<113> vss vdd vss wl<113> / cell_PIM
XI25242 vss vss in1<115> in2<115> vss vdd vss wl<115> / cell_PIM
XI25241 vss vss in1<117> in2<117> vss vdd vss wl<117> / cell_PIM
XI25240 vss vss in1<116> in2<116> vss vdd vss wl<116> / cell_PIM
XI25239 vss vss in1<118> in2<118> vss vdd vss wl<118> / cell_PIM
XI25243 vss vss in1<114> in2<114> vss vdd vss wl<114> / cell_PIM
XI25237 vss vss in1<122> in2<122> vss vdd vss wl<122> / cell_PIM
XI25236 vss vss in1<121> in2<121> vss vdd vss wl<121> / cell_PIM
XI25235 vss vss in1<120> in2<120> vss vdd vss wl<120> / cell_PIM
XI25234 vss vss in1<123> in2<123> vss vdd vss wl<123> / cell_PIM
XI25238 vss vss in1<119> in2<119> vss vdd vss wl<119> / cell_PIM
XI25232 vss vss in1<127> in2<127> vss vdd vss wl<127> / cell_PIM
XI25231 vss vss in1<126> in2<126> vss vdd vss wl<126> / cell_PIM
XI25230 vss vss in1<125> in2<125> vss vdd vss wl<125> / cell_PIM
XI25229 vss vss in1<124> in2<124> vss vdd vss wl<124> / cell_PIM
XI25233 vss vss vdd vdd vss vdd vss vss / cell_PIM
XI25228 vss vss vdd vdd vss vdd vss vss / cell_PIM2
XI25227 vss vss in1<0> in2<0> vss vdd vss wl<0> / cell_PIM2
XI25226 vss vss in1<1> in2<1> vss vdd vss wl<1> / cell_PIM2
XI25225 vss vss in1<2> in2<2> vss vdd vss wl<2> / cell_PIM2
XI25224 vss vss in1<4> in2<4> vss vdd vss wl<4> / cell_PIM2
XI25222 vss vss in1<5> in2<5> vss vdd vss wl<5> / cell_PIM2
XI25221 vss vss in1<6> in2<6> vss vdd vss wl<6> / cell_PIM2
XI25220 vss vss in1<7> in2<7> vss vdd vss wl<7> / cell_PIM2
XI25219 vss vss in1<8> in2<8> vss vdd vss wl<8> / cell_PIM2
XI25223 vss vss in1<3> in2<3> vss vdd vss wl<3> / cell_PIM2
XI25217 vss vss in1<10> in2<10> vss vdd vss wl<10> / cell_PIM2
XI25216 vss vss in1<11> in2<11> vss vdd vss wl<11> / cell_PIM2
XI25215 vss vss in1<12> in2<12> vss vdd vss wl<12> / cell_PIM2
XI25214 vss vss in1<13> in2<13> vss vdd vss wl<13> / cell_PIM2
XI25218 vss vss in1<9> in2<9> vss vdd vss wl<9> / cell_PIM2
XI25212 vss vss in1<15> in2<15> vss vdd vss wl<15> / cell_PIM2
XI25211 vss vss in1<16> in2<16> vss vdd vss wl<16> / cell_PIM2
XI25210 vss vss in1<17> in2<17> vss vdd vss wl<17> / cell_PIM2
XI25209 vss vss in1<18> in2<18> vss vdd vss wl<18> / cell_PIM2
XI25213 vss vss in1<14> in2<14> vss vdd vss wl<14> / cell_PIM2
XI25208 vss vss in1<19> in2<19> vss vdd vss wl<19> / cell_PIM2
XI25207 vss vss in1<20> in2<20> vss vdd vss wl<20> / cell_PIM2
XI25206 vss vss in1<21> in2<21> vss vdd vss wl<21> / cell_PIM2
XI25205 vss vss in1<22> in2<22> vss vdd vss wl<22> / cell_PIM2
XI25204 vss vss in1<23> in2<23> vss vdd vss wl<23> / cell_PIM2
XI25202 vss vss in1<25> in2<25> vss vdd vss wl<25> / cell_PIM2
XI25201 vss vss in1<26> in2<26> vss vdd vss wl<26> / cell_PIM2
XI25200 vss vss in1<27> in2<27> vss vdd vss wl<27> / cell_PIM2
XI25199 vss vss in1<28> in2<28> vss vdd vss wl<28> / cell_PIM2
XI25203 vss vss in1<24> in2<24> vss vdd vss wl<24> / cell_PIM2
XI25197 vss vss in1<30> in2<30> vss vdd vss wl<30> / cell_PIM2
XI25196 vss vss in1<31> in2<31> vss vdd vss wl<31> / cell_PIM2
XI25195 vss vss in1<32> in2<32> vss vdd vss wl<32> / cell_PIM2
XI25194 vss vss in1<33> in2<33> vss vdd vss wl<33> / cell_PIM2
XI25198 vss vss in1<29> in2<29> vss vdd vss wl<29> / cell_PIM2
XI25192 vss vss in1<35> in2<35> vss vdd vss wl<35> / cell_PIM2
XI25191 vss vss in1<36> in2<36> vss vdd vss wl<36> / cell_PIM2
XI25190 vss vss in1<37> in2<37> vss vdd vss wl<37> / cell_PIM2
XI25189 vss vss in1<38> in2<38> vss vdd vss wl<38> / cell_PIM2
XI25193 vss vss in1<34> in2<34> vss vdd vss wl<34> / cell_PIM2
XI25188 vss vss in1<39> in2<39> vss vdd vss wl<39> / cell_PIM2
XI25187 vss vss in1<40> in2<40> vss vdd vss wl<40> / cell_PIM2
XI25186 vss vss in1<41> in2<41> vss vdd vss wl<41> / cell_PIM2
XI25185 vss vss in1<42> in2<42> vss vdd vss wl<42> / cell_PIM2
XI25184 vss vss in1<43> in2<43> vss vdd vss wl<43> / cell_PIM2
XI25182 vss vss in1<45> in2<45> vss vdd vss wl<45> / cell_PIM2
XI25181 vss vss in1<46> in2<46> vss vdd vss wl<46> / cell_PIM2
XI25180 vss vss in1<47> in2<47> vss vdd vss wl<47> / cell_PIM2
XI25179 vss vss in1<48> in2<48> vss vdd vss wl<48> / cell_PIM2
XI25183 vss vss in1<44> in2<44> vss vdd vss wl<44> / cell_PIM2
XI25177 vss vss in1<50> in2<50> vss vdd vss wl<50> / cell_PIM2
XI25176 vss vss in1<51> in2<51> vss vdd vss wl<51> / cell_PIM2
XI25175 vss vss in1<52> in2<52> vss vdd vss wl<52> / cell_PIM2
XI25174 vss vss in1<53> in2<53> vss vdd vss wl<53> / cell_PIM2
XI25178 vss vss in1<49> in2<49> vss vdd vss wl<49> / cell_PIM2
XI25172 vss vss in1<55> in2<55> vss vdd vss wl<55> / cell_PIM2
XI25171 vss vss in1<56> in2<56> vss vdd vss wl<56> / cell_PIM2
XI25170 vss vss in1<57> in2<57> vss vdd vss wl<57> / cell_PIM2
XI25169 vss vss in1<58> in2<58> vss vdd vss wl<58> / cell_PIM2
XI25173 vss vss in1<54> in2<54> vss vdd vss wl<54> / cell_PIM2
XI25168 vss vss in1<59> in2<59> vss vdd vss wl<59> / cell_PIM2
XI25167 vss vss in1<60> in2<60> vss vdd vss wl<60> / cell_PIM2
XI25166 vss vss in1<61> in2<61> vss vdd vss wl<61> / cell_PIM2
XI25165 vss vss in1<62> in2<62> vss vdd vss wl<62> / cell_PIM2
XI25164 vss vss in1<63> in2<63> vss vdd vss wl<63> / cell_PIM2
XI25162 vss vss in1<65> in2<65> vss vdd vss wl<65> / cell_PIM2
XI25161 vss vss in1<66> in2<66> vss vdd vss wl<66> / cell_PIM2
XI25160 vss vss in1<67> in2<67> vss vdd vss wl<67> / cell_PIM2
XI25159 vss vss in1<68> in2<68> vss vdd vss wl<68> / cell_PIM2
XI25163 vss vss in1<64> in2<64> vss vdd vss wl<64> / cell_PIM2
XI25157 vss vss in1<70> in2<70> vss vdd vss wl<70> / cell_PIM2
XI25156 vss vss in1<71> in2<71> vss vdd vss wl<71> / cell_PIM2
XI25155 vss vss in1<72> in2<72> vss vdd vss wl<72> / cell_PIM2
XI25154 vss vss in1<73> in2<73> vss vdd vss wl<73> / cell_PIM2
XI25158 vss vss in1<69> in2<69> vss vdd vss wl<69> / cell_PIM2
XI25152 vss vss in1<75> in2<75> vss vdd vss wl<75> / cell_PIM2
XI25151 vss vss in1<76> in2<76> vss vdd vss wl<76> / cell_PIM2
XI25150 vss vss in1<77> in2<77> vss vdd vss wl<77> / cell_PIM2
XI25149 vss vss in1<78> in2<78> vss vdd vss wl<78> / cell_PIM2
XI25153 vss vss in1<74> in2<74> vss vdd vss wl<74> / cell_PIM2
XI25148 vss vss in1<79> in2<79> vss vdd vss wl<79> / cell_PIM2
XI25147 vss vss in1<80> in2<80> vss vdd vss wl<80> / cell_PIM2
XI25146 vss vss in1<81> in2<81> vss vdd vss wl<81> / cell_PIM2
XI25145 vss vss in1<82> in2<82> vss vdd vss wl<82> / cell_PIM2
XI25144 vss vss in1<83> in2<83> vss vdd vss wl<83> / cell_PIM2
XI25142 vss vss in1<85> in2<85> vss vdd vss wl<85> / cell_PIM2
XI25141 vss vss in1<86> in2<86> vss vdd vss wl<86> / cell_PIM2
XI25140 vss vss in1<87> in2<87> vss vdd vss wl<87> / cell_PIM2
XI25139 vss vss in1<88> in2<88> vss vdd vss wl<88> / cell_PIM2
XI25143 vss vss in1<84> in2<84> vss vdd vss wl<84> / cell_PIM2
XI25137 vss vss in1<90> in2<90> vss vdd vss wl<90> / cell_PIM2
XI25136 vss vss in1<91> in2<91> vss vdd vss wl<91> / cell_PIM2
XI25135 vss vss in1<92> in2<92> vss vdd vss wl<92> / cell_PIM2
XI25134 vss vss in1<93> in2<93> vss vdd vss wl<93> / cell_PIM2
XI25138 vss vss in1<89> in2<89> vss vdd vss wl<89> / cell_PIM2
XI25132 vss vss in1<95> in2<95> vss vdd vss wl<95> / cell_PIM2
XI25131 vss vss in1<96> in2<96> vss vdd vss wl<96> / cell_PIM2
XI25130 vss vss in1<97> in2<97> vss vdd vss wl<97> / cell_PIM2
XI25129 vss vss in1<98> in2<98> vss vdd vss wl<98> / cell_PIM2
XI25133 vss vss in1<94> in2<94> vss vdd vss wl<94> / cell_PIM2
XI25128 vss vss in1<99> in2<99> vss vdd vss wl<99> / cell_PIM2
XI25127 vss vss in1<100> in2<100> vss vdd vss wl<100> / cell_PIM2
XI25126 vss vss in1<101> in2<101> vss vdd vss wl<101> / cell_PIM2
XI25125 vss vss in1<102> in2<102> vss vdd vss wl<102> / cell_PIM2
XI25124 vss vss in1<103> in2<103> vss vdd vss wl<103> / cell_PIM2
XI25122 vss vss in1<105> in2<105> vss vdd vss wl<105> / cell_PIM2
XI25121 vss vss in1<106> in2<106> vss vdd vss wl<106> / cell_PIM2
XI25120 vss vss in1<107> in2<107> vss vdd vss wl<107> / cell_PIM2
XI25119 vss vss in1<108> in2<108> vss vdd vss wl<108> / cell_PIM2
XI25123 vss vss in1<104> in2<104> vss vdd vss wl<104> / cell_PIM2
XI25117 vss vss in1<110> in2<110> vss vdd vss wl<110> / cell_PIM2
XI25116 vss vss in1<111> in2<111> vss vdd vss wl<111> / cell_PIM2
XI25115 vss vss in1<112> in2<112> vss vdd vss wl<112> / cell_PIM2
XI25114 vss vss in1<113> in2<113> vss vdd vss wl<113> / cell_PIM2
XI25118 vss vss in1<109> in2<109> vss vdd vss wl<109> / cell_PIM2
XI25112 vss vss in1<115> in2<115> vss vdd vss wl<115> / cell_PIM2
XI25111 vss vss in1<116> in2<116> vss vdd vss wl<116> / cell_PIM2
XI25110 vss vss in1<117> in2<117> vss vdd vss wl<117> / cell_PIM2
XI25109 vss vss in1<118> in2<118> vss vdd vss wl<118> / cell_PIM2
XI25113 vss vss in1<114> in2<114> vss vdd vss wl<114> / cell_PIM2
XI25108 vss vss in1<119> in2<119> vss vdd vss wl<119> / cell_PIM2
XI25107 vss vss in1<120> in2<120> vss vdd vss wl<120> / cell_PIM2
XI25106 vss vss in1<121> in2<121> vss vdd vss wl<121> / cell_PIM2
XI25105 vss vss in1<122> in2<122> vss vdd vss wl<122> / cell_PIM2
XI25104 vss vss in1<123> in2<123> vss vdd vss wl<123> / cell_PIM2
XI25102 vss vss in1<127> in2<127> vss vdd vss wl<127> / cell_PIM2
XI25101 vss vss in1<126> in2<126> vss vdd vss wl<126> / cell_PIM2
XI25100 vss vss in1<125> in2<125> vss vdd vss wl<125> / cell_PIM2
XI25099 vss vss in1<124> in2<124> vss vdd vss wl<124> / cell_PIM2
XI25103 vss vss vdd vdd vss vdd vss vss / cell_PIM2
XI33745 bl<0> bl<1> bl<2> bl<3> cbl<0> cbl<1> col_en in1<0> in1<1> in1<2> 
+ in1<4> in1<3> in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> 
+ in1<13> in1<14> in1<15> in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> 
+ in1<22> in1<23> in1<24> in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> 
+ in1<31> in1<32> in1<33> in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> 
+ in1<40> in1<41> in1<42> in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> 
+ in1<49> in1<50> in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> 
+ in1<58> in1<59> in1<60> in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> 
+ in1<67> in1<68> in1<69> in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> 
+ in1<76> in1<77> in1<78> in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> 
+ in1<85> in1<86> in1<87> in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> 
+ in1<94> in1<95> in1<96> in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> 
+ in1<103> in1<104> in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> 
+ in1<111> in1<112> in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> 
+ in1<119> in1<120> in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> 
+ in1<127> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> 
+ in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> 
+ in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> 
+ in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> 
+ in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> 
+ in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> 
+ in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> 
+ in2<63> in2<64> in2<65> in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> 
+ in2<72> in2<73> in2<74> in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> 
+ in2<81> in2<82> in2<83> in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> 
+ in2<90> in2<91> in2<92> in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> 
+ in2<99> in2<100> in2<101> in2<102> in2<103> in2<104> in2<105> in2<106> 
+ in2<107> in2<108> in2<109> in2<110> in2<111> in2<112> in2<113> in2<114> 
+ in2<115> in2<116> in2<117> in2<118> in2<119> in2<120> in2<121> in2<122> 
+ in2<123> in2<124> in2<125> in2<126> in2<127> reg_en sel<0> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> 
+ wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> wl<20> 
+ wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> 
+ wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> wl<42> 
+ wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> wl<53> 
+ wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> wl<64> 
+ wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> wl<75> 
+ wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> wl<86> 
+ wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> wl<97> 
+ wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127> / array_test_cel_2
XI33751 bl<12> bl<13> bl<14> bl<15> cbl<6> cbl<7> col_en in1<0> in1<1> in1<2> 
+ in1<4> in1<3> in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> 
+ in1<13> in1<14> in1<15> in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> 
+ in1<22> in1<23> in1<24> in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> 
+ in1<31> in1<32> in1<33> in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> 
+ in1<40> in1<41> in1<42> in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> 
+ in1<49> in1<50> in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> 
+ in1<58> in1<59> in1<60> in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> 
+ in1<67> in1<68> in1<69> in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> 
+ in1<76> in1<77> in1<78> in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> 
+ in1<85> in1<86> in1<87> in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> 
+ in1<94> in1<95> in1<96> in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> 
+ in1<103> in1<104> in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> 
+ in1<111> in1<112> in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> 
+ in1<119> in1<120> in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> 
+ in1<127> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> 
+ in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> 
+ in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> 
+ in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> 
+ in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> 
+ in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> 
+ in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> 
+ in2<63> in2<64> in2<65> in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> 
+ in2<72> in2<73> in2<74> in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> 
+ in2<81> in2<82> in2<83> in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> 
+ in2<90> in2<91> in2<92> in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> 
+ in2<99> in2<100> in2<101> in2<102> in2<103> in2<104> in2<105> in2<106> 
+ in2<107> in2<108> in2<109> in2<110> in2<111> in2<112> in2<113> in2<114> 
+ in2<115> in2<116> in2<117> in2<118> in2<119> in2<120> in2<121> in2<122> 
+ in2<123> in2<124> in2<125> in2<126> in2<127> reg_en sel<3> sl<12> sl<13> 
+ sl<14> sl<15> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> 
+ wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> 
+ wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> 
+ wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> 
+ wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> 
+ wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> 
+ wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> 
+ wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> 
+ wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> 
+ wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127> / array_test_cel_2
XI33749 bl<4> bl<5> bl<6> bl<7> cbl<2> cbl<3> col_en in1<0> in1<1> in1<2> 
+ in1<4> in1<3> in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> 
+ in1<13> in1<14> in1<15> in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> 
+ in1<22> in1<23> in1<24> in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> 
+ in1<31> in1<32> in1<33> in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> 
+ in1<40> in1<41> in1<42> in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> 
+ in1<49> in1<50> in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> 
+ in1<58> in1<59> in1<60> in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> 
+ in1<67> in1<68> in1<69> in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> 
+ in1<76> in1<77> in1<78> in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> 
+ in1<85> in1<86> in1<87> in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> 
+ in1<94> in1<95> in1<96> in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> 
+ in1<103> in1<104> in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> 
+ in1<111> in1<112> in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> 
+ in1<119> in1<120> in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> 
+ in1<127> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> 
+ in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> 
+ in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> 
+ in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> 
+ in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> 
+ in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> 
+ in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> 
+ in2<63> in2<64> in2<65> in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> 
+ in2<72> in2<73> in2<74> in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> 
+ in2<81> in2<82> in2<83> in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> 
+ in2<90> in2<91> in2<92> in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> 
+ in2<99> in2<100> in2<101> in2<102> in2<103> in2<104> in2<105> in2<106> 
+ in2<107> in2<108> in2<109> in2<110> in2<111> in2<112> in2<113> in2<114> 
+ in2<115> in2<116> in2<117> in2<118> in2<119> in2<120> in2<121> in2<122> 
+ in2<123> in2<124> in2<125> in2<126> in2<127> reg_en sel<1> sl<4> sl<5> sl<6> 
+ sl<7> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> 
+ wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> wl<20> 
+ wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> 
+ wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> wl<42> 
+ wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> wl<53> 
+ wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> wl<64> 
+ wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> wl<75> 
+ wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> wl<86> 
+ wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> wl<97> 
+ wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127> / array_test_cel_2
XI33750 bl<8> bl<9> bl<10> bl<11> cbl<4> cbl<5> col_en in1<0> in1<1> in1<2> 
+ in1<4> in1<3> in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> 
+ in1<13> in1<14> in1<15> in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> 
+ in1<22> in1<23> in1<24> in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> 
+ in1<31> in1<32> in1<33> in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> 
+ in1<40> in1<41> in1<42> in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> 
+ in1<49> in1<50> in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> 
+ in1<58> in1<59> in1<60> in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> 
+ in1<67> in1<68> in1<69> in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> 
+ in1<76> in1<77> in1<78> in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> 
+ in1<85> in1<86> in1<87> in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> 
+ in1<94> in1<95> in1<96> in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> 
+ in1<103> in1<104> in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> 
+ in1<111> in1<112> in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> 
+ in1<119> in1<120> in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> 
+ in1<127> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> 
+ in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> 
+ in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> 
+ in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> 
+ in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> 
+ in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> 
+ in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> 
+ in2<63> in2<64> in2<65> in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> 
+ in2<72> in2<73> in2<74> in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> 
+ in2<81> in2<82> in2<83> in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> 
+ in2<90> in2<91> in2<92> in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> 
+ in2<99> in2<100> in2<101> in2<102> in2<103> in2<104> in2<105> in2<106> 
+ in2<107> in2<108> in2<109> in2<110> in2<111> in2<112> in2<113> in2<114> 
+ in2<115> in2<116> in2<117> in2<118> in2<119> in2<120> in2<121> in2<122> 
+ in2<123> in2<124> in2<125> in2<126> in2<127> reg_en sel<2> sl<8> sl<9> 
+ sl<10> sl<11> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> 
+ wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> 
+ wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> 
+ wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> 
+ wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> 
+ wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> 
+ wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> 
+ wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> 
+ wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> 
+ wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127> / array_test_cel_2
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    Dtriger
* View Name:    schematic
************************************************************************

.SUBCKT Dtriger cp d q qn rdn sdn vdd vss
*.PININFO cp:I d:I rdn:I sdn:I q:O qn:O vdd:B vss:B
XI12 vdd vss net10 sdn net19 net27 / 3nand
XI9 vdd vss rdn net27 cp net19 / 3nand
XI8 vdd vss qn net19 sdn q / 3nand
XI11 vdd vss net18 rdn d net10 / 3nand
XI6 vdd vss rdn net18 q qn / 3nand
XI10 vdd vss cp net10 net19 net18 / 3nand
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor IN0 IN1 OUT VDD VSS
*.PININFO IN0:B IN1:B OUT:B VDD:B VSS:B
XNM2 OUT IN1 VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM3 OUT IN0 VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XPM3 OUT IN1 net018 VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM0 net018 IN0 VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    Tgate2
* View Name:    schematic
************************************************************************

.SUBCKT Tgate2 IN OE OEN OUT VDD VSS
*.PININFO IN:B OE:B OEN:B OUT:B VDD:B VSS:B
XNM2 OUT OE IN VSS n12ll_mis_ckt MR=1 L=80n W=600n
XPM0 IN OEN OUT VDD p12ll_mis_ckt MR=1 L=80n W=600n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    countercell
* View Name:    schematic
************************************************************************

.SUBCKT countercell col_en cp q<0> q<1> q<2> q<3> q<4> q<5> setn vdd vss
*.PININFO col_en:I cp:I setn:I q<0>:O q<1>:O q<2>:O q<3>:O q<4>:O q<5>:O vdd:B 
*.PININFO vss:B
XI34 net050 net052 net053 net052 setn vdd vdd vss / Dtriger
XI28 net046 net048 net049 net048 setn vdd vdd vss / Dtriger
XI29 net048 net050 net051 net050 setn vdd vdd vss / Dtriger
XI23 net61 net046 net047 net046 setn vdd vdd vss / Dtriger
XI8 net59 net61 net62 net61 setn vdd vdd vss / Dtriger
XI0 clk net59 net60 net59 setn vdd vdd vss / Dtriger
XI41 clk_en clk_en_n vdd vss / inv1
XI5 col_en col_en_n vdd vss / inv1
XI31 net056 q<4> vdd vss / inv1
XI25 net058 q<2> vdd vss / inv1
XI18 net76 q<1> vdd vss / inv1
XI17 net77 q<0> vdd vss / inv1
XI30 net051 net056 vdd vss / inv1
XI33 net053 net055 vdd vss / inv1
XI32 net055 q<5> vdd vss / inv1
XI26 net057 q<3> vdd vss / inv1
XI27 net049 net057 vdd vss / inv1
XI24 net047 net058 vdd vss / inv1
XI3 net60 net77 vdd vss / inv1
XI7 net62 net76 vdd vss / inv1
XI38 vdd vss q<5> q<4> q<3> and_1 / 3nand
XI37 vdd vss q<2> q<1> q<0> and_0 / 3nand
XI40 and_1 and_0 net018 vdd vss / nor
XI39 col_en_n and_0 net019 vdd vss / nor
XI22 net019 net018 clk_en vdd vss / nor
XI10 cp clk_en clk_en_n clk vdd vss / Tgate2
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    countercell2
* View Name:    schematic
************************************************************************

.SUBCKT countercell2 adco<0> adco<1> col_en q<0> q<1> q<2> q<3> q<4> q<5> q<6> 
+ q<7> q<8> q<9> q<10> q<11> setn vdd vss
*.PININFO adco<0>:I adco<1>:I col_en:I setn:I q<0>:O q<1>:O q<2>:O q<3>:O 
*.PININFO q<4>:O q<5>:O q<6>:O q<7>:O q<8>:O q<9>:O q<10>:O q<11>:O vdd:B vss:B
XI1 col_en adco<1> q<6> q<7> q<8> q<9> q<10> q<11> setn vdd vss / countercell
XI0 col_en adco<0> q<0> q<1> q<2> q<3> q<4> q<5> setn vdd vss / countercell
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    counter
* View Name:    schematic
************************************************************************

.SUBCKT counter adc<0> adc<1> adc<2> adc<3> adc<4> adc<5> adc<6> adc<7> adc<8> 
+ adc<9> adc<10> adc<11> adc<12> adc<13> adc<14> adc<15> adc<16> adc<17> 
+ adc<18> adc<19> adc<20> adc<21> adc<22> adc<23> adc<24> adc<25> adc<26> 
+ adc<27> adc<28> adc<29> adc<30> adc<31> col_en d<0> d<1> d<2> d<3> d<4> d<5> 
+ d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> d<16> d<17> d<18> 
+ d<19> d<20> d<21> d<22> d<23> d<24> d<25> d<26> d<27> d<28> d<29> d<30> 
+ d<31> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> 
+ q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> 
+ q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> 
+ q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> 
+ q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> 
+ q<61> q<62> q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> 
+ q<73> q<74> q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> 
+ q<85> q<86> q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> 
+ q<97> q<98> q<99> q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> 
+ q<108> q<109> q<110> q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> 
+ q<119> q<120> q<121> q<122> q<123> q<124> q<125> q<126> q<127> q<128> q<129> 
+ q<130> q<131> q<132> q<133> q<134> q<135> q<136> q<137> q<138> q<139> q<140> 
+ q<141> q<142> q<143> q<144> q<145> q<146> q<147> q<148> q<149> q<150> q<151> 
+ q<152> q<153> q<154> q<155> q<156> q<157> q<158> q<159> q<160> q<161> q<162> 
+ q<163> q<164> q<165> q<166> q<167> q<168> q<169> q<170> q<171> q<172> q<173> 
+ q<174> q<175> q<176> q<177> q<178> q<179> q<180> q<181> q<182> q<183> q<184> 
+ q<185> q<186> q<187> q<188> q<189> q<190> q<191> set vdd vss
*.PININFO adc<0>:I adc<1>:I adc<2>:I adc<3>:I adc<4>:I adc<5>:I adc<6>:I 
*.PININFO adc<7>:I adc<8>:I adc<9>:I adc<10>:I adc<11>:I adc<12>:I adc<13>:I 
*.PININFO adc<14>:I adc<15>:I adc<16>:I adc<17>:I adc<18>:I adc<19>:I 
*.PININFO adc<20>:I adc<21>:I adc<22>:I adc<23>:I adc<24>:I adc<25>:I 
*.PININFO adc<26>:I adc<27>:I adc<28>:I adc<29>:I adc<30>:I adc<31>:I col_en:I 
*.PININFO set:I q<0>:O q<1>:O q<2>:O q<3>:O q<4>:O q<5>:O q<6>:O q<7>:O q<8>:O 
*.PININFO q<9>:O q<10>:O q<11>:O q<12>:O q<13>:O q<14>:O q<15>:O q<16>:O 
*.PININFO q<17>:O q<18>:O q<19>:O q<20>:O q<21>:O q<22>:O q<23>:O q<24>:O 
*.PININFO q<25>:O q<26>:O q<27>:O q<28>:O q<29>:O q<30>:O q<31>:O q<32>:O 
*.PININFO q<33>:O q<34>:O q<35>:O q<36>:O q<37>:O q<38>:O q<39>:O q<40>:O 
*.PININFO q<41>:O q<42>:O q<43>:O q<44>:O q<45>:O q<46>:O q<47>:O q<48>:O 
*.PININFO q<49>:O q<50>:O q<51>:O q<52>:O q<53>:O q<54>:O q<55>:O q<56>:O 
*.PININFO q<57>:O q<58>:O q<59>:O q<60>:O q<61>:O q<62>:O q<63>:O q<64>:O 
*.PININFO q<65>:O q<66>:O q<67>:O q<68>:O q<69>:O q<70>:O q<71>:O q<72>:O 
*.PININFO q<73>:O q<74>:O q<75>:O q<76>:O q<77>:O q<78>:O q<79>:O q<80>:O 
*.PININFO q<81>:O q<82>:O q<83>:O q<84>:O q<85>:O q<86>:O q<87>:O q<88>:O 
*.PININFO q<89>:O q<90>:O q<91>:O q<92>:O q<93>:O q<94>:O q<95>:O q<96>:O 
*.PININFO q<97>:O q<98>:O q<99>:O q<100>:O q<101>:O q<102>:O q<103>:O q<104>:O 
*.PININFO q<105>:O q<106>:O q<107>:O q<108>:O q<109>:O q<110>:O q<111>:O 
*.PININFO q<112>:O q<113>:O q<114>:O q<115>:O q<116>:O q<117>:O q<118>:O 
*.PININFO q<119>:O q<120>:O q<121>:O q<122>:O q<123>:O q<124>:O q<125>:O 
*.PININFO q<126>:O q<127>:O q<128>:O q<129>:O q<130>:O q<131>:O q<132>:O 
*.PININFO q<133>:O q<134>:O q<135>:O q<136>:O q<137>:O q<138>:O q<139>:O 
*.PININFO q<140>:O q<141>:O q<142>:O q<143>:O q<144>:O q<145>:O q<146>:O 
*.PININFO q<147>:O q<148>:O q<149>:O q<150>:O q<151>:O q<152>:O q<153>:O 
*.PININFO q<154>:O q<155>:O q<156>:O q<157>:O q<158>:O q<159>:O q<160>:O 
*.PININFO q<161>:O q<162>:O q<163>:O q<164>:O q<165>:O q<166>:O q<167>:O 
*.PININFO q<168>:O q<169>:O q<170>:O q<171>:O q<172>:O q<173>:O q<174>:O 
*.PININFO q<175>:O q<176>:O q<177>:O q<178>:O q<179>:O q<180>:O q<181>:O 
*.PININFO q<182>:O q<183>:O q<184>:O q<185>:O q<186>:O q<187>:O q<188>:O 
*.PININFO q<189>:O q<190>:O q<191>:O d<0>:B d<1>:B d<2>:B d<3>:B d<4>:B d<5>:B 
*.PININFO d<6>:B d<7>:B d<8>:B d<9>:B d<10>:B d<11>:B d<12>:B d<13>:B d<14>:B 
*.PININFO d<15>:B d<16>:B d<17>:B d<18>:B d<19>:B d<20>:B d<21>:B d<22>:B 
*.PININFO d<23>:B d<24>:B d<25>:B d<26>:B d<27>:B d<28>:B d<29>:B d<30>:B 
*.PININFO d<31>:B vdd:B vss:B
XI2 adc<0> adc<1> col_en q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> 
+ q<10> q<11> setn vdd vss / countercell2
XI20 set setn vdd vss / inv4
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv2
* View Name:    schematic
************************************************************************

.SUBCKT inv2 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=60n W=900n
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=60n W=1.8u
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv8
* View Name:    schematic
************************************************************************

.SUBCKT inv8 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=1u
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=1u
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    master
* View Name:    schematic
************************************************************************

.SUBCKT master a<0> a<1> a<2> a<3> a<4> a<5> a<6> a<7> a_col<0> a_col<1> 
+ a_row<0> a_row<1> a_row<2> a_row<3> a_row<4> a_row<5> a_row<6> clk comp 
+ en_acc_col en_acc_row entime inbit model model_ set set_ set_comp time<0> 
+ time<1> time<2> time<3> vdd vss wait wrt wrt_ wrtbuf_
*.PININFO a<0>:I a<1>:I a<2>:I a<3>:I a<4>:I a<5>:I a<6>:I a<7>:I clk:I comp:I 
*.PININFO inbit:I model:I set:I wait:I wrt:I a_col<0>:O a_col<1>:O a_row<0>:O 
*.PININFO a_row<1>:O a_row<2>:O a_row<3>:O a_row<4>:O a_row<5>:O a_row<6>:O 
*.PININFO en_acc_col:O en_acc_row:O entime:O model_:O set_:O set_comp:O 
*.PININFO time<0>:O time<1>:O time<2>:O time<3>:O wrt_:O wrtbuf_:O vdd:B vss:B
XI102 net015 waitb vdd vss / inv2
XI114 net018 net049 vdd vss / inv2
XI113 net019 net018 vdd vss / inv2
XI116 net0100 net039 vdd vss / inv2
XI115 net016 net0100 vdd vss / inv2
XI122 net0101 ab<8> vdd vss / inv2
XI46 net077 net074 vdd vss / inv2
XI1<0> net094<0> ab<0> vdd vss / inv2
XI1<1> net094<1> ab<1> vdd vss / inv2
XI1<2> net094<2> ab<2> vdd vss / inv2
XI1<3> net094<3> ab<3> vdd vss / inv2
XI1<4> net094<4> ab<4> vdd vss / inv2
XI1<5> net094<5> ab<5> vdd vss / inv2
XI1<6> net094<6> ab<6> vdd vss / inv2
XI1<7> net094<7> ab<7> vdd vss / inv2
XI7 net051 compb vdd vss / inv2
XI5 net050 setb vdd vss / inv2
XI13 net040 readb vdd vss / inv2
XI15 net039 inbitb vdd vss / inv2
XI2 net049 modelb vdd vss / inv2
XI17 net038 wrtbufb vdd vss / inv2
XI11 net053 wrtb vdd vss / inv2
XI101 wait net015 vdd vss / inv8
XI0<0> a<0> net094<0> vdd vss / inv8
XI0<1> a<1> net094<1> vdd vss / inv8
XI0<2> a<2> net094<2> vdd vss / inv8
XI0<3> a<3> net094<3> vdd vss / inv8
XI0<4> a<4> net094<4> vdd vss / inv8
XI0<5> a<5> net094<5> vdd vss / inv8
XI0<6> a<6> net094<6> vdd vss / inv8
XI0<7> a<7> net094<7> vdd vss / inv8
XI65<0> net084<0> a_row<0> vdd vss / inv8
XI65<1> net084<1> a_row<1> vdd vss / inv8
XI65<2> net084<2> a_row<2> vdd vss / inv8
XI65<3> net084<3> a_row<3> vdd vss / inv8
XI65<4> net084<4> a_row<4> vdd vss / inv8
XI65<5> net084<5> a_row<5> vdd vss / inv8
XI65<6> net084<6> a_row<6> vdd vss / inv8
XI70<0> net085<0> a_col<0> vdd vss / inv8
XI70<1> net085<1> a_col<1> vdd vss / inv8
XI72<0> net059<0> a_read<0> vdd vss / inv8
XI72<1> net059<1> a_read<1> vdd vss / inv8
XI72<2> net059<2> a_read<2> vdd vss / inv8
XI72<3> net059<3> a_read<3> vdd vss / inv8
XI68<0> net060<0> a_inbuf<0> vdd vss / inv8
XI68<1> net060<1> a_inbuf<1> vdd vss / inv8
XI68<2> net060<2> a_inbuf<2> vdd vss / inv8
XI68<3> net060<3> a_inbuf<3> vdd vss / inv8
XI68<4> net060<4> a_inbuf<4> vdd vss / inv8
XI59 net064 eninbuf vdd vss / inv8
XI58 net067 en_acc_col vdd vss / inv8
XI56 net068 en_acc_row vdd vss / inv8
XI53 net069 enread vdd vss / inv8
XI49 net070 set_comp vdd vss / inv8
XI43 net076 clk_write vdd vss / inv8
XI39 net062 clk_read vdd vss / inv8
XI31 net080 set_ vdd vss / inv8
XI30 net081 model_ vdd vss / inv8
XI8 clk net052 vdd vss / inv8
XI9 net052 clkb vdd vss / inv8
XI6 comp net051 vdd vss / inv8
XI4 set net050 vdd vss / inv8
XI14 inbit net016 vdd vss / inv8
XI12 vss net040 vdd vss / inv8
XI16 vss net038 vdd vss / inv8
XI26 net061 wrtbuf_ vdd vss / inv8
XI19 net06 wrt_ vdd vss / inv8
XI3 model net019 vdd vss / inv8
XI123 vss net0101 vdd vss / inv8
XI10 wrt net053 vdd vss / inv8
XI112 clkcharge net026 net022 vdd vss / nand
XI110 clkcharge net025 net023 vdd vss / nand
XI108 clkcharge net027 net024 vdd vss / nand
XI106 clkcharge net029 net028 vdd vss / nand
XI104 clkb net012 net097 vdd vss / nand
XI99 net0126 inbitb net0132 vdd vss / nand
XI96 compb modelb net0128 vdd vss / nand
XI93 net066 inbitn net065 vdd vss / nand
XI90 compb modelb net0122 vdd vss / nand
XI87 net0137 inbitb net0124 vdd vss / nand
XI84 compb modeln net0121 vdd vss / nand
XI81 net0131 inbitn net0120 vdd vss / nand
XI78 compb modeln net0136 vdd vss / nand
XI47 net074 clkb net075 vdd vss / nand
XI37 clkb readb net079 vdd vss / nand
XI20 clkb wrtbufb net014 vdd vss / nand
XI18 clkb wrtb net013 vdd vss / nand
XI111 net022 time<0> vdd vss / inv4
XI109 net023 time<1> vdd vss / inv4
XI107 net024 time<2> vdd vss / inv4
XI105 net028 time<3> vdd vss / inv4
XI103 net097 clkcharge vdd vss / inv4
XI98 net0132 net029 vdd vss / inv4
XI97 net0128 net0126 vdd vss / inv4
XI92 net065 net027 vdd vss / inv4
XI91 net0122 net066 vdd vss / inv4
XI86 net0124 net025 vdd vss / inv4
XI85 net0121 net0137 vdd vss / inv4
XI69<0> ab<7> net085<0> vdd vss / inv4
XI69<1> ab<8> net085<1> vdd vss / inv4
XI75 inbitb inbitn vdd vss / inv4
XI67<0> ab<0> net060<0> vdd vss / inv4
XI67<1> ab<1> net060<1> vdd vss / inv4
XI67<2> ab<2> net060<2> vdd vss / inv4
XI67<3> ab<3> net060<3> vdd vss / inv4
XI67<4> ab<4> net060<4> vdd vss / inv4
XI71<0> ab<0> net059<0> vdd vss / inv4
XI71<1> ab<1> net059<1> vdd vss / inv4
XI71<2> ab<2> net059<2> vdd vss / inv4
XI71<3> ab<3> net059<3> vdd vss / inv4
XI80 net0120 net026 vdd vss / inv4
XI79 net0136 net0131 vdd vss / inv4
XI66<0> ab<0> net084<0> vdd vss / inv4
XI66<1> ab<1> net084<1> vdd vss / inv4
XI66<2> ab<2> net084<2> vdd vss / inv4
XI66<3> ab<3> net084<3> vdd vss / inv4
XI66<4> ab<4> net084<4> vdd vss / inv4
XI66<5> ab<5> net084<5> vdd vss / inv4
XI66<6> ab<6> net084<6> vdd vss / inv4
XI119 net095 net012 vdd vss / inv4
XI60 net061 net064 vdd vss / inv4
XI57 net06 net067 vdd vss / inv4
XI55 net06 net068 vdd vss / inv4
XI54 net062 net069 vdd vss / inv4
XI52 net072 entime vdd vss / inv4
XI50 entime net070 vdd vss / inv4
XI48 net075 net073 vdd vss / inv4
XI44 net073 net076 vdd vss / inv4
XI38 net079 net078 vdd vss / inv4
XI40 net078 net062 vdd vss / inv4
XI82 modelb modeln vdd vss / inv4
XI32 setb net080 vdd vss / inv4
XI29 modelb net081 vdd vss / inv4
XI25 net011 net06 vdd vss / inv4
XI28 net082 net061 vdd vss / inv4
XI27 net014 net082 vdd vss / inv4
XI22 net013 net011 vdd vss / inv4
XI118 waitb setb net095 vdd vss / nor
XI51 setb compb net072 vdd vss / nor
XI45 wrtb wrtbufb net077 vdd vss / nor
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    SA
* View Name:    schematic
************************************************************************

.SUBCKT SA in1 in2 out vb vdd vss
*.PININFO in1:I in2:I vb:I out:B vdd:B vss:B
XPM2 net021 in2 net16 vdd p12ll_mis_ckt MR=1 L=120n W=600n
XPM3 net019 in1 net16 vdd p12ll_mis_ckt MR=1 L=120n W=600n
XPM0 net07 net07 vdd vdd p12ll_mis_ckt MR=1 L=120n W=2.4u
XPM1 net16 vb vdd vdd p12ll_mis_ckt MR=1 L=120n W=600n
XPM4 out net07 vdd vdd p12ll_mis_ckt MR=1 L=120n W=19.2u
XNM1 net07 net019 vss vss n12ll_mis_ckt MR=1 L=120n W=1.2u
XNM2 net021 net019 vss vss n12ll_mis_ckt MR=1 L=120n W=300n
XNM3 out net021 vss vss n12ll_mis_ckt MR=1 L=87n W=9.6u
XNM0 net019 net019 vss vss n12ll_mis_ckt MR=1 L=120n W=300n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    bias
* View Name:    schematic
************************************************************************

.SUBCKT bias set set_comp vb vb2 vb3 vdd vss
*.PININFO set:I set_comp:I vb:O vb2:O vb3:O vdd:B vss:B
XI36 net010 setn setb vb vdd vss / Tgate
XI38 vb2 setb setn net09 vdd vss / Tgate
XI37 net018 setb setn vb vdd vss / Tgate
XI39 vbr set_compb set_compn net010 vdd vss / Tgate
XI35 setn setb vdd vss / inv4
XI34 set setn vdd vss / inv4
XI10 set_compn set_compb vdd vss / inv4
XI9 set_comp set_compn vdd vss / inv4
XI25 vb net010 net018 net09 vdd vss / SA
XPM0 vbr vbr vdd vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM2 vb3 set_compn net05 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM6 vb3 set_compn net027 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM7 vb2 set_compn net011 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM9 vb2 set_compn net028 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM10 net09 setb vdd vdd p12ll_mis_ckt MR=1 L=600n W=600n
XPM1 vbr vbr vdd vdd p12ll_mis_ckt MR=1 L=600n W=1u
XNM6 vbr set_compb net026 vss n12ll_mis_ckt MR=1 L=600n W=1u
XNM15 vb2 vb2 vss vss n12ll_mis_ckt MR=1 L=600n W=500n
XNM16 vbr set_compb net1 vss n12ll_mis_ckt MR=1 L=600n W=1u
XNM10 vb3 vb3 vss vss n12ll_mis_ckt MR=1 L=600n W=600n
XNM12 vb2 vb2 vss vss n12ll_mis_ckt MR=1 L=600n W=500n
XNM11 vb3 vb3 vss vss n12ll_mis_ckt MR=1 L=600n W=600n
XR7 vdd net028 rhrpo_ckt M=1 W=2u L=800u
XR0 net026 vss rhrpo_ckt M=1 W=2u L=10u
XR1 net1 vss rhrpo_ckt M=1 W=2u L=10u
XR6 vdd net011 rhrpo_ckt M=1 W=2u L=800u
XR9 vdd net027 rhrpo_ckt M=1 W=2u L=80u
XR8 vdd net05 rhrpo_ckt M=1 W=2u L=80u
XC8 vb2 vss mom_2t_ckt LF=5u NF=10 TM=3 BM=1 MR=1
XC9 vb vss mom_2t_ckt LF=5u NF=20 TM=3 BM=1 MR=1
XC5 vb3 vss mom_2t_ckt LF=5u NF=10 TM=3 BM=1 MR=1
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv0_5
* View Name:    schematic
************************************************************************

.SUBCKT inv0_5 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    invz
* View Name:    schematic
************************************************************************

.SUBCKT invz IN OE OEN OUT VDD VSS
*.PININFO IN:B OE:B OEN:B OUT:B VDD:B VSS:B
XPM3 OUT OEN net13 VDD p12ll_mis_ckt MR=1 L=80n W=200n
XPM2 net13 IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XNM3 net14 IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
XNM2 OUT OE net14 VSS n12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv0_3
* View Name:    schematic
************************************************************************

.SUBCKT inv0_3 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    SA2
* View Name:    schematic
************************************************************************

.SUBCKT SA2 in1 in2 out vb vdd vss
*.PININFO in1:I in2:I vb:I vdd:I vss:I out:B
XNM8 net015 net015 vss vss n12ll_mis_ckt MR=1 L=80n W=150n
XNM0 net01 net015 vss vss n12ll_mis_ckt MR=1 L=80n W=150n
XNM7 net07 net015 vss vss n12ll_mis_ckt MR=1 L=80n W=300n
XNM9 out net01 vss vss n12ll_mis_ckt MR=1 L=80n W=300n
XPM7 net07 net07 vdd vdd p12ll_mis_ckt MR=1 L=80n W=600n
XPM5 net01 in2 net26 vdd p12ll_mis_ckt MR=1 L=80n W=300n
XPM4 net26 vb vdd vdd p12ll_mis_ckt MR=1 L=80n W=300n
XPM8 net015 in1 net26 vdd p12ll_mis_ckt MR=1 L=80n W=300n
XPM9 out net07 vdd vdd p12ll_mis_ckt MR=1 L=80n W=600n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    ADCcell_2
* View Name:    schematic
************************************************************************

.SUBCKT ADCcell_2 cbl model set set_comp set_compn setn vb vb2 vb3 vdd vss x<5>
*.PININFO cbl:I model:I set:I set_comp:I set_compn:I setn:I vb:I vb2:I vb3:I 
*.PININFO vdd:I vss:I x<5>:O
XI23 net54 net014 vdd vss / inv0_5
XI22 x<1> set net54 vdd vss / nor
XNM5 Vc x<3> vss vss n12ll_mis_ckt MR=1 L=80n W=1.2u
XNM4 vss set_compn x<1> vss n12ll_mis_ckt MR=1 L=80n W=300n
XNM3 net016 bc Vc vss n12ll_mis_ckt MR=1 L=80n W=1.2u
XNM2 cbl vb3 net016 vss n12ll_mis_ckt MR=1 L=80n W=600n
XNM6 Vc set vss vss n12ll_mis_ckt MR=1 L=80n W=600n
XI7 x<0> set_comp set_compn x<1> vdd vss / invz
XI1 cbl set setn vb vdd vss / Tgate
XI3<0> x<1> x<2> vdd vss / inv0_3
XI3<1> x<2> x<3> vdd vss / inv0_3
XI3<2> x<3> x<4> vdd vss / inv0_3
XI10 Vc model_n model net013 vdd vss / Tgate2
XI8 x<4> x<5> vdd vss / inv1
XI11 model model_n vdd vss / inv1
XI5 net014 bc vdd vss / inv1
XI0 Vc vb x<0> vb2 vdd vss / SA2
XC2 cbl vss mom_2t_ckt LF=20u NF=32 TM=3 BM=1 MR=1
XC5 Vc vss mom_2t_ckt LF=1u NF=6 TM=3 BM=1 MR=1
XC6 net013 vss mom_2t_ckt LF=1u NF=24 TM=3 BM=1 MR=1
XPM0 vdd set_comp vb2 vdd p12ll_mis_ckt MR=1 L=80n W=1.2u
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    ADC
* View Name:    schematic
************************************************************************

.SUBCKT ADC adc<0> adc<1> adc<2> adc<3> adc<4> adc<5> adc<6> adc<7> adc<8> 
+ adc<9> adc<10> adc<11> adc<12> adc<13> adc<14> adc<15> adc<16> adc<17> 
+ adc<18> adc<19> adc<20> adc<21> adc<22> adc<23> adc<24> adc<25> adc<26> 
+ adc<27> adc<28> adc<29> adc<30> adc<31> cbl<0> cbl<1> cbl<2> cbl<3> cbl<4> 
+ cbl<5> cbl<6> cbl<7> cbl<8> cbl<9> cbl<10> cbl<11> cbl<12> cbl<13> cbl<14> 
+ cbl<15> cbl<16> cbl<17> cbl<18> cbl<19> cbl<20> cbl<21> cbl<22> cbl<23> 
+ cbl<24> cbl<25> cbl<26> cbl<27> cbl<28> cbl<29> cbl<30> cbl<31> d<0> d<1> 
+ d<2> d<3> d<4> d<5> d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> 
+ d<16> d<17> d<18> d<19> d<20> d<21> d<22> d<23> d<24> d<25> d<26> d<27> 
+ d<28> d<29> d<30> d<31> model set set_comp vdd vss
*.PININFO cbl<0>:I cbl<1>:I cbl<2>:I cbl<3>:I cbl<4>:I cbl<5>:I cbl<6>:I 
*.PININFO cbl<7>:I cbl<8>:I cbl<9>:I cbl<10>:I cbl<11>:I cbl<12>:I cbl<13>:I 
*.PININFO cbl<14>:I cbl<15>:I cbl<16>:I cbl<17>:I cbl<18>:I cbl<19>:I 
*.PININFO cbl<20>:I cbl<21>:I cbl<22>:I cbl<23>:I cbl<24>:I cbl<25>:I 
*.PININFO cbl<26>:I cbl<27>:I cbl<28>:I cbl<29>:I cbl<30>:I cbl<31>:I model:I 
*.PININFO set:I set_comp:I adc<0>:O adc<1>:O adc<2>:O adc<3>:O adc<4>:O 
*.PININFO adc<5>:O adc<6>:O adc<7>:O adc<8>:O adc<9>:O adc<10>:O adc<11>:O 
*.PININFO adc<12>:O adc<13>:O adc<14>:O adc<15>:O adc<16>:O adc<17>:O 
*.PININFO adc<18>:O adc<19>:O adc<20>:O adc<21>:O adc<22>:O adc<23>:O 
*.PININFO adc<24>:O adc<25>:O adc<26>:O adc<27>:O adc<28>:O adc<29>:O 
*.PININFO adc<30>:O adc<31>:O d<0>:B d<1>:B d<2>:B d<3>:B d<4>:B d<5>:B d<6>:B 
*.PININFO d<7>:B d<8>:B d<9>:B d<10>:B d<11>:B d<12>:B d<13>:B d<14>:B d<15>:B 
*.PININFO d<16>:B d<17>:B d<18>:B d<19>:B d<20>:B d<21>:B d<22>:B d<23>:B 
*.PININFO d<24>:B d<25>:B d<26>:B d<27>:B d<28>:B d<29>:B d<30>:B d<31>:B 
*.PININFO vdd:B vss:B
XI7 set_compn set_compb vdd vss / inv4
XI6 set_comp set_compn vdd vss / inv4
XI3 modelbn modelb vdd vss / inv4
XI2 model modelbn vdd vss / inv4
XI1 setbn setb vdd vss / inv4
XI16 set setbn vdd vss / inv4
XI5 setb set_compb vb vb2 vb3 vdd vss / bias
XI41 cbl<0> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<0> / 
+ ADCcell_2
XI15 cbl<4> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<4> / 
+ ADCcell_2
XI14 cbl<6> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<6> / 
+ ADCcell_2
XI13 cbl<7> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<7> / 
+ ADCcell_2
XI12 cbl<5> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<5> / 
+ ADCcell_2
XI11 cbl<2> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<2> / 
+ ADCcell_2
XI10 cbl<3> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<3> / 
+ ADCcell_2
XI9 cbl<1> modelb setb set_compb set_compn setbn vb vb2 vb3 vdd vss adc<1> / 
+ ADCcell_2
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Writecell_2
* View Name:    schematic
************************************************************************

.SUBCKT Writecell_2 VDD VSS bl<0> bl<1> col<0> col<1> d reg_en sl<0> sl<1> wrt 
+ wrtbuf
*.PININFO col<0>:I col<1>:I d:I reg_en:I wrt:I wrtbuf:I bl<0>:O bl<1>:O 
*.PININFO sl<0>:O sl<1>:O VDD:B VSS:B
XI26 wrt reg_en net021 VDD VSS / nor
XI15 wrt_regen wrtbuf net013 VDD VSS / nor
XI12 wrtalln d wdnb VDD VSS / nor
XI5 wrtalln dn wdns VDD VSS / nor
XI25 net021 wrt_regen VDD VSS / inv2
XI13 wdnb wdps VDD VSS / inv2
XI6 wdns wdpb VDD VSS / inv2
XI7 d dn VDD VSS / inv2
XI3<0> wrt_regen col<0> net017<0> VDD VSS / nand
XI3<1> wrt_regen col<1> net017<1> VDD VSS / nand
XI9<0> bl<0> net018<0> net019<0> tBL VDD VSS / Tgate
XI9<1> bl<1> net018<1> net019<1> tBL VDD VSS / Tgate
XI10<0> sl<0> net018<0> net019<0> tSL VDD VSS / Tgate
XI10<1> sl<1> net018<1> net019<1> tSL VDD VSS / Tgate
XI16 net013 wrtall VDD VSS / inv1
XI11 wrtall wrtalln VDD VSS / inv1
XI14<0> net017<0> net018<0> VDD VSS / inv1
XI14<1> net017<1> net018<1> VDD VSS / inv1
XI8<0> net018<0> net019<0> VDD VSS / inv1
XI8<1> net018<1> net019<1> VDD VSS / inv1
XPM2 tBL wdpb VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM1 tSL wdps VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XNM0 tBL wdnb VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM1 tSL wdns VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Writedriver
* View Name:    schematic
************************************************************************

.SUBCKT Writedriver bl<0> bl<1> bl<2> bl<3> bl<4> bl<5> bl<6> bl<7> bl<8> 
+ bl<9> bl<10> bl<11> bl<12> bl<13> bl<14> bl<15> bl<16> bl<17> bl<18> bl<19> 
+ bl<20> bl<21> bl<22> bl<23> bl<24> bl<25> bl<26> bl<27> bl<28> bl<29> bl<30> 
+ bl<31> bl<32> bl<33> bl<34> bl<35> bl<36> bl<37> bl<38> bl<39> bl<40> bl<41> 
+ bl<42> bl<43> bl<44> bl<45> bl<46> bl<47> bl<48> bl<49> bl<50> bl<51> bl<52> 
+ bl<53> bl<54> bl<55> bl<56> bl<57> bl<58> bl<59> bl<60> bl<61> bl<62> bl<63> 
+ cbl<0> cbl<1> cbl<2> cbl<3> cbl<4> cbl<5> cbl<6> cbl<7> cbl<8> cbl<9> 
+ cbl<10> cbl<11> cbl<12> cbl<13> cbl<14> cbl<15> cbl<16> cbl<17> cbl<18> 
+ cbl<19> cbl<20> cbl<21> cbl<22> cbl<23> cbl<24> cbl<25> cbl<26> cbl<27> 
+ cbl<28> cbl<29> cbl<30> cbl<31> col<0> col<1> d<0> d<1> d<2> d<3> d<4> d<5> 
+ d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> d<16> d<17> d<18> 
+ d<19> d<20> d<21> d<22> d<23> d<24> d<25> d<26> d<27> d<28> d<29> d<30> 
+ d<31> reg_en sl<0> sl<1> sl<2> sl<3> sl<4> sl<5> sl<6> sl<7> sl<8> sl<9> 
+ sl<10> sl<11> sl<12> sl<13> sl<14> sl<15> sl<16> sl<17> sl<18> sl<19> sl<20> 
+ sl<21> sl<22> sl<23> sl<24> sl<25> sl<26> sl<27> sl<28> sl<29> sl<30> sl<31> 
+ sl<32> sl<33> sl<34> sl<35> sl<36> sl<37> sl<38> sl<39> sl<40> sl<41> sl<42> 
+ sl<43> sl<44> sl<45> sl<46> sl<47> sl<48> sl<49> sl<50> sl<51> sl<52> sl<53> 
+ sl<54> sl<55> sl<56> sl<57> sl<58> sl<59> sl<60> sl<61> sl<62> sl<63> vdd 
+ vss wrt wrtbuf
*.PININFO col<0>:I col<1>:I d<0>:I d<1>:I d<2>:I d<3>:I d<4>:I d<5>:I d<6>:I 
*.PININFO d<7>:I d<8>:I d<9>:I d<10>:I d<11>:I d<12>:I d<13>:I d<14>:I d<15>:I 
*.PININFO d<16>:I d<17>:I d<18>:I d<19>:I d<20>:I d<21>:I d<22>:I d<23>:I 
*.PININFO d<24>:I d<25>:I d<26>:I d<27>:I d<28>:I d<29>:I d<30>:I d<31>:I 
*.PININFO reg_en:I wrt:I wrtbuf:I bl<0>:O bl<1>:O bl<2>:O bl<3>:O bl<4>:O 
*.PININFO bl<5>:O bl<6>:O bl<7>:O bl<8>:O bl<9>:O bl<10>:O bl<11>:O bl<12>:O 
*.PININFO bl<13>:O bl<14>:O bl<15>:O bl<16>:O bl<17>:O bl<18>:O bl<19>:O 
*.PININFO bl<20>:O bl<21>:O bl<22>:O bl<23>:O bl<24>:O bl<25>:O bl<26>:O 
*.PININFO bl<27>:O bl<28>:O bl<29>:O bl<30>:O bl<31>:O bl<32>:O bl<33>:O 
*.PININFO bl<34>:O bl<35>:O bl<36>:O bl<37>:O bl<38>:O bl<39>:O bl<40>:O 
*.PININFO bl<41>:O bl<42>:O bl<43>:O bl<44>:O bl<45>:O bl<46>:O bl<47>:O 
*.PININFO bl<48>:O bl<49>:O bl<50>:O bl<51>:O bl<52>:O bl<53>:O bl<54>:O 
*.PININFO bl<55>:O bl<56>:O bl<57>:O bl<58>:O bl<59>:O bl<60>:O bl<61>:O 
*.PININFO bl<62>:O bl<63>:O sl<0>:O sl<1>:O sl<2>:O sl<3>:O sl<4>:O sl<5>:O 
*.PININFO sl<6>:O sl<7>:O sl<8>:O sl<9>:O sl<10>:O sl<11>:O sl<12>:O sl<13>:O 
*.PININFO sl<14>:O sl<15>:O sl<16>:O sl<17>:O sl<18>:O sl<19>:O sl<20>:O 
*.PININFO sl<21>:O sl<22>:O sl<23>:O sl<24>:O sl<25>:O sl<26>:O sl<27>:O 
*.PININFO sl<28>:O sl<29>:O sl<30>:O sl<31>:O sl<32>:O sl<33>:O sl<34>:O 
*.PININFO sl<35>:O sl<36>:O sl<37>:O sl<38>:O sl<39>:O sl<40>:O sl<41>:O 
*.PININFO sl<42>:O sl<43>:O sl<44>:O sl<45>:O sl<46>:O sl<47>:O sl<48>:O 
*.PININFO sl<49>:O sl<50>:O sl<51>:O sl<52>:O sl<53>:O sl<54>:O sl<55>:O 
*.PININFO sl<56>:O sl<57>:O sl<58>:O sl<59>:O sl<60>:O sl<61>:O sl<62>:O 
*.PININFO sl<63>:O cbl<0>:B cbl<1>:B cbl<2>:B cbl<3>:B cbl<4>:B cbl<5>:B 
*.PININFO cbl<6>:B cbl<7>:B cbl<8>:B cbl<9>:B cbl<10>:B cbl<11>:B cbl<12>:B 
*.PININFO cbl<13>:B cbl<14>:B cbl<15>:B cbl<16>:B cbl<17>:B cbl<18>:B 
*.PININFO cbl<19>:B cbl<20>:B cbl<21>:B cbl<22>:B cbl<23>:B cbl<24>:B 
*.PININFO cbl<25>:B cbl<26>:B cbl<27>:B cbl<28>:B cbl<29>:B cbl<30>:B 
*.PININFO cbl<31>:B vdd:B vss:B
XI50 vdd vss bl<31> bl<63> col<0> col<1> d<31> reg_en sl<31> sl<63> wrt wrtbuf 
+ / Writecell_2
XI49 vdd vss bl<30> bl<62> col<0> col<1> d<30> reg_en sl<30> sl<62> wrt wrtbuf 
+ / Writecell_2
XI48 vdd vss bl<29> bl<61> col<0> col<1> d<29> reg_en sl<29> sl<61> wrt wrtbuf 
+ / Writecell_2
XI47 vdd vss bl<28> bl<60> col<0> col<1> d<28> reg_en sl<28> sl<60> wrt wrtbuf 
+ / Writecell_2
XI46 vdd vss bl<27> bl<59> col<0> col<1> d<27> reg_en sl<27> sl<59> wrt wrtbuf 
+ / Writecell_2
XI45 vdd vss bl<26> bl<58> col<0> col<1> d<26> reg_en sl<26> sl<58> wrt wrtbuf 
+ / Writecell_2
XI44 vdd vss bl<25> bl<57> col<0> col<1> d<25> reg_en sl<25> sl<57> wrt wrtbuf 
+ / Writecell_2
XI43 vdd vss bl<24> bl<56> col<0> col<1> d<24> reg_en sl<24> sl<56> wrt wrtbuf 
+ / Writecell_2
XI42 vdd vss bl<23> bl<55> col<0> col<1> d<23> reg_en sl<23> sl<55> wrt wrtbuf 
+ / Writecell_2
XI41 vdd vss bl<22> bl<54> col<0> col<1> d<22> reg_en sl<22> sl<54> wrt wrtbuf 
+ / Writecell_2
XI40 vdd vss bl<21> bl<53> col<0> col<1> d<21> reg_en sl<21> sl<53> wrt wrtbuf 
+ / Writecell_2
XI39 vdd vss bl<20> bl<52> col<0> col<1> d<20> reg_en sl<20> sl<52> wrt wrtbuf 
+ / Writecell_2
XI38 vdd vss bl<19> bl<51> col<0> col<1> d<19> reg_en sl<19> sl<51> wrt wrtbuf 
+ / Writecell_2
XI37 vdd vss bl<18> bl<50> col<0> col<1> d<18> reg_en sl<18> sl<50> wrt wrtbuf 
+ / Writecell_2
XI36 vdd vss bl<17> bl<49> col<0> col<1> d<17> reg_en sl<17> sl<49> wrt wrtbuf 
+ / Writecell_2
XI35 vdd vss bl<16> bl<48> col<0> col<1> d<16> reg_en sl<16> sl<48> wrt wrtbuf 
+ / Writecell_2
XI16 vdd vss bl<15> bl<47> col<0> col<1> d<15> reg_en sl<15> sl<47> wrt wrtbuf 
+ / Writecell_2
XI15 vdd vss bl<14> bl<46> col<0> col<1> d<14> reg_en sl<14> sl<46> wrt wrtbuf 
+ / Writecell_2
XI14 vdd vss bl<13> bl<45> col<0> col<1> d<13> reg_en sl<13> sl<45> wrt wrtbuf 
+ / Writecell_2
XI13 vdd vss bl<12> bl<44> col<0> col<1> d<12> reg_en sl<12> sl<44> wrt wrtbuf 
+ / Writecell_2
XI12 vdd vss bl<11> bl<43> col<0> col<1> d<11> reg_en sl<11> sl<43> wrt wrtbuf 
+ / Writecell_2
XI11 vdd vss bl<10> bl<42> col<0> col<1> d<10> reg_en sl<10> sl<42> wrt wrtbuf 
+ / Writecell_2
XI10 vdd vss bl<9> bl<41> col<0> col<1> d<9> reg_en sl<9> sl<41> wrt wrtbuf / 
+ Writecell_2
XI9 vdd vss bl<8> bl<40> col<0> col<1> d<8> reg_en sl<8> sl<40> wrt wrtbuf / 
+ Writecell_2
XI8 vdd vss bl<7> bl<39> col<0> col<1> d<7> reg_en sl<7> sl<39> wrt wrtbuf / 
+ Writecell_2
XI7 vdd vss bl<6> bl<38> col<0> col<1> d<6> reg_en sl<6> sl<38> wrt wrtbuf / 
+ Writecell_2
XI6 vdd vss bl<5> bl<37> col<0> col<1> d<5> reg_en sl<5> sl<37> wrt wrtbuf / 
+ Writecell_2
XI5 vdd vss bl<4> bl<36> col<0> col<1> d<4> reg_en sl<4> sl<36> wrt wrtbuf / 
+ Writecell_2
XI4 vdd vss bl<3> bl<35> col<0> col<1> d<3> reg_en sl<3> sl<35> wrt wrtbuf / 
+ Writecell_2
XI3 vdd vss bl<2> bl<34> col<0> col<1> d<2> reg_en sl<2> sl<34> wrt wrtbuf / 
+ Writecell_2
XI2 vdd vss bl<1> bl<33> col<0> col<1> d<1> reg_en sl<1> sl<33> wrt wrtbuf / 
+ Writecell_2
XI1 vdd vss bl<0> bl<32> col<0> col<1> d<0> reg_en sl<0> sl<32> wrt wrtbuf / 
+ Writecell_2
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    3x8decoder
* View Name:    schematic
************************************************************************

.SUBCKT 3x8decoder in<0> in<1> in<2> out<0> out<1> out<2> out<3> out<4> out<5> 
+ out<6> out<7> vdd vss
*.PININFO in<0>:I in<1>:I in<2>:I out<0>:O out<1>:O out<2>:O out<3>:O out<4>:O 
*.PININFO out<5>:O out<6>:O out<7>:O vdd:B vss:B
XI1 vdd vss inn<2> in<0> in<1> out<4> out<5> out<6> out<7> / 2x4decoder
XI0 vdd vss in<2> in<0> in<1> out<0> out<1> out<2> out<3> / 2x4decoder
XI2 in<2> inn<2> vdd vss / inv1
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    4x16decoder
* View Name:    schematic
************************************************************************

.SUBCKT 4x16decoder VDD VSS en in<0> in<1> in<2> in<3> out<0> out<1> out<2> 
+ out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11> out<12> 
+ out<13> out<14> out<15>
*.PININFO en:I in<0>:I in<1>:I in<2>:I in<3>:I out<0>:O out<1>:O out<2>:O 
*.PININFO out<3>:O out<4>:O out<5>:O out<6>:O out<7>:O out<8>:O out<9>:O 
*.PININFO out<10>:O out<11>:O out<12>:O out<13>:O out<14>:O out<15>:O VDD:B 
*.PININFO VSS:B
XI15 VDD VSS en in<2> in<3> b<0> b<1> b<2> b<3> / 2x4decoder
XI0 VDD VSS en in<0> in<1> c<0> c<1> c<2> c<3> / 2x4decoder
XI73 net173 out<15> VDD VSS / inv4
XI70 net174 out<14> VDD VSS / inv4
XI69 net175 out<13> VDD VSS / inv4
XI67 net176 out<12> VDD VSS / inv4
XI81 net092 out<11> VDD VSS / inv4
XI78 net097 out<10> VDD VSS / inv4
XI77 net179 out<9> VDD VSS / inv4
XI75 net180 out<8> VDD VSS / inv4
XI65 net0112 out<7> VDD VSS / inv4
XI62 net182 out<6> VDD VSS / inv4
XI61 net183 out<5> VDD VSS / inv4
XI59 net0127 out<4> VDD VSS / inv4
XI57 net185 out<3> VDD VSS / inv4
XI54 net0137 out<2> VDD VSS / inv4
XI53 net187 out<1> VDD VSS / inv4
XI51 net188 out<0> VDD VSS / inv4
XI8 c<2> b<2> net097 VDD VSS / nand
XI7 c<3> b<2> net092 VDD VSS / nand
XI6 c<3> b<1> net0112 VDD VSS / nand
XI5 c<2> b<1> net182 VDD VSS / nand
XI4 c<0> b<1> net0127 VDD VSS / nand
XI3 c<1> b<1> net183 VDD VSS / nand
XI2 c<3> b<0> net185 VDD VSS / nand
XI1 c<2> b<0> net0137 VDD VSS / nand
XI9 c<0> b<2> net180 VDD VSS / nand
XI10 c<1> b<2> net179 VDD VSS / nand
XI11 c<1> b<3> net175 VDD VSS / nand
XI12 c<0> b<3> net176 VDD VSS / nand
XI13 c<2> b<3> net174 VDD VSS / nand
XI14 c<3> b<3> net173 VDD VSS / nand
XI50 c<0> b<0> net188 VDD VSS / nand
XI52 c<1> b<0> net187 VDD VSS / nand
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    access_decoder
* View Name:    schematic
************************************************************************

.SUBCKT access_decoder a_col<0> a_col<1> a_row<0> a_row<1> a_row<2> a_row<3> 
+ a_row<4> a_row<5> a_row<6> col<0> col<1> en_acc_col en_acc_row group<0> 
+ group<1> group<2> group<3> group<4> group<5> group<6> group<7> reg_en 
+ row16<0> row16<1> row16<2> row16<3> row16<4> row16<5> row16<6> row16<7> 
+ row16<8> row16<9> row16<10> row16<11> row16<12> row16<13> row16<14> 
+ row16<15> vdd vss wrt wrtbuf
*.PININFO a_col<0>:I a_col<1>:I a_row<0>:I a_row<1>:I a_row<2>:I a_row<3>:I 
*.PININFO a_row<4>:I a_row<5>:I a_row<6>:I en_acc_col:I en_acc_row:I reg_en:I 
*.PININFO col<0>:O col<1>:O group<0>:O group<1>:O group<2>:O group<3>:O 
*.PININFO group<4>:O group<5>:O group<6>:O group<7>:O row16<0>:O row16<1>:O 
*.PININFO row16<2>:O row16<3>:O row16<4>:O row16<5>:O row16<6>:O row16<7>:O 
*.PININFO row16<8>:O row16<9>:O row16<10>:O row16<11>:O row16<12>:O 
*.PININFO row16<13>:O row16<14>:O row16<15>:O vdd:B vss:B wrt:B wrtbuf:B
XI0 a_row<0> a_row<1> a_row<2> group<0> group<1> group<2> group<3> group<4> 
+ group<5> group<6> group<7> vdd vss / 3x8decoder
XI1 vdd vss en_acc_row a_row<3> a_row<4> a_row<5> a_row<6> row16<0> row16<1> 
+ row16<2> row16<3> row16<4> row16<5> row16<6> row16<7> row16<8> row16<9> 
+ row16<10> row16<11> row16<12> row16<13> row16<14> row16<15> / 4x16decoder
XI2 vdd vss en_acc_col_decode a_col<0> a_col<1> col<0> col<1> net2 net1 / 
+ 2x4decoder
XI23 en_acc_col_n reg_en en_acc_col_decode VDD VSS / nor
XI24 en_acc_col en_acc_col_n VDD VSS / inv2
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    delaycell_editable
* View Name:    schematic
************************************************************************

.SUBCKT delaycell_editable VDD VSS in out
*.PININFO in:I out:O VDD:B VSS:B
XI1<0> x<0> x<1> VDD VSS / inv0_3
XI1<1> x<1> x<2> VDD VSS / inv0_3
XI1<2> x<2> x<3> VDD VSS / inv0_3
XI1<3> x<3> x<4> VDD VSS / inv0_3
XI1<4> x<4> x<5> VDD VSS / inv0_3
XI1<5> x<5> x<6> VDD VSS / inv0_3
XI1<6> x<6> x<7> VDD VSS / inv0_3
XI1<7> x<7> x<8> VDD VSS / inv0_3
XI1<8> x<8> x<9> VDD VSS / inv0_3
XI1<9> x<9> x<10> VDD VSS / inv0_3
XI0 in x<0> VDD VSS / inv0_3
XI2 x<10> out VDD VSS / inv1
XPM4 out x<10> out VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM2 x<0> in x<0> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<0> x<1> x<0> x<1> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<1> x<2> x<1> x<2> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<2> x<3> x<2> x<3> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<3> x<4> x<3> x<4> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<4> x<5> x<4> x<5> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<5> x<6> x<5> x<6> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<6> x<7> x<6> x<7> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<7> x<8> x<7> x<8> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<8> x<9> x<8> x<9> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<9> x<10> x<9> x<10> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XNM6 out x<10> out VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<0> x<1> x<0> x<1> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<1> x<2> x<1> x<2> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<2> x<3> x<2> x<3> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<3> x<4> x<3> x<4> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<4> x<5> x<4> x<5> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<5> x<6> x<5> x<6> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<6> x<7> x<6> x<7> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<7> x<8> x<7> x<8> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<8> x<9> x<8> x<9> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<9> x<10> x<9> x<10> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM0 x<0> in x<0> VSS n12ll_mis_ckt MR=1 L=80n W=400n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate entime in1 in2 q<0> q<1> q<2> q<3> time<0> time<1> time<2> 
+ time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I time<0>:I time<1>:I time<2>:I 
*.PININFO time<3>:I in1:O in2:O vdd:B vss:B
XI21 net014 net013 net025 vdd vss / nor
XI17 net15 net14 net19 vdd vss / nor
XI12 net19 net011 net18 vdd vss / nor
XI22 net024 net026 vdd vss / inv4
XI13 net027 net17 vdd vss / inv4
XI23 net026 in2 vdd vss / inv8
XI14 net17 in1 vdd vss / inv8
XI20 net013 net014 net027 vdd vss / nand
XI7 q<3> time<3> net10 vdd vss / nand
XI6 q<2> time<2> net11 vdd vss / nand
XI16 net11 net10 net14 vdd vss / nand
XI3 q<1> time<1> net12 vdd vss / nand
XI15 net13 net12 net15 vdd vss / nand
XI0 q<0> time<0> net13 vdd vss / nand
XI24 net025 net024 vdd vss / inv1
XI19 net18 net013 vdd vss / inv1
XI30 entime net011 vdd vss / inv1
XI27 vdd vss net013 net014 / delaycell_editable
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_2
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_2 entime in1<0> in1<1> in2<0> in2<1> q<0> q<1> q<2> 
+ q<3> q<4> q<5> q<6> q<7> time<0> time<1> time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO time<0>:I time<1>:I time<2>:I time<3>:I in1<0>:O in1<1>:O in2<0>:O 
*.PININFO in2<1>:O vdd:B vss:B
XI0 entime in1<0> in2<0> q<0> q<1> q<2> q<3> time<0> time<1> time<2> time<3> 
+ vdd vss / Tgenerate
XI1 entime in1<1> in2<1> q<4> q<5> q<6> q<7> time<0> time<1> time<2> time<3> 
+ vdd vss / Tgenerate
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_4
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_4 entime in1<0> in1<1> in1<2> in1<3> in2<0> in2<1> 
+ in2<2> in2<3> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> 
+ q<12> q<13> q<14> q<15> time<0> time<1> time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO time<0>:I time<1>:I time<2>:I time<3>:I in1<0>:O in1<1>:O in1<2>:O 
*.PININFO in1<3>:O in2<0>:O in2<1>:O in2<2>:O in2<3>:O vdd:B vss:B
XI128 entime in1<0> in1<1> in2<0> in2<1> q<0> q<1> q<2> q<3> q<4> q<5> q<6> 
+ q<7> time<0> time<1> time<2> time<3> vdd vss / Tgenerate_array_2
XI129 entime in1<2> in1<3> in2<2> in2<3> q<8> q<9> q<10> q<11> q<12> q<13> 
+ q<14> q<15> time<0> time<1> time<2> time<3> vdd vss / Tgenerate_array_2
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_8
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_8 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> 
+ in1<6> in1<7> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> q<0> 
+ q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> 
+ q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> 
+ q<27> q<28> q<29> q<30> q<31> time<0> time<1> time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO q<16>:I q<17>:I q<18>:I q<19>:I q<20>:I q<21>:I q<22>:I q<23>:I 
*.PININFO q<24>:I q<25>:I q<26>:I q<27>:I q<28>:I q<29>:I q<30>:I q<31>:I 
*.PININFO time<0>:I time<1>:I time<2>:I time<3>:I in1<0>:O in1<1>:O in1<2>:O 
*.PININFO in1<3>:O in1<4>:O in1<5>:O in1<6>:O in1<7>:O in2<0>:O in2<1>:O 
*.PININFO in2<2>:O in2<3>:O in2<4>:O in2<5>:O in2<6>:O in2<7>:O vdd:B vss:B
XI130 entimeb in1<0> in1<1> in1<2> in1<3> in2<0> in2<1> in2<2> in2<3> q<0> 
+ q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> 
+ q<15> timeb<0> timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate_array_4
XI131 entimeb in1<4> in1<5> in1<6> in1<7> in2<4> in2<5> in2<6> in2<7> q<16> 
+ q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> q<27> q<28> 
+ q<29> q<30> q<31> timeb<0> timeb<1> timeb<2> timeb<3> vdd vss / 
+ Tgenerate_array_4
XI3 entime net09 vdd vss / inv4
XI25<0> time<0> net011<0> vdd vss / inv4
XI25<1> time<1> net011<1> vdd vss / inv4
XI25<2> time<2> net011<2> vdd vss / inv4
XI25<3> time<3> net011<3> vdd vss / inv4
XI2 net09 entimeb vdd vss / inv8
XI1<0> net011<0> timeb<0> vdd vss / inv8
XI1<1> net011<1> timeb<1> vdd vss / inv8
XI1<2> net011<2> timeb<2> vdd vss / inv8
XI1<3> net011<3> timeb<3> vdd vss / inv8
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_16
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_16 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> 
+ in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> 
+ in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> 
+ in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> q<0> q<1> q<2> q<3> q<4> 
+ q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> q<15> q<16> q<17> 
+ q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> q<27> q<28> q<29> 
+ q<30> q<31> q<32> q<33> q<34> q<35> q<36> q<37> q<38> q<39> q<40> q<41> 
+ q<42> q<43> q<44> q<45> q<46> q<47> q<48> q<49> q<50> q<51> q<52> q<53> 
+ q<54> q<55> q<56> q<57> q<58> q<59> q<60> q<61> q<62> q<63> time<0> time<1> 
+ time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO q<16>:I q<17>:I q<18>:I q<19>:I q<20>:I q<21>:I q<22>:I q<23>:I 
*.PININFO q<24>:I q<25>:I q<26>:I q<27>:I q<28>:I q<29>:I q<30>:I q<31>:I 
*.PININFO q<32>:I q<33>:I q<34>:I q<35>:I q<36>:I q<37>:I q<38>:I q<39>:I 
*.PININFO q<40>:I q<41>:I q<42>:I q<43>:I q<44>:I q<45>:I q<46>:I q<47>:I 
*.PININFO q<48>:I q<49>:I q<50>:I q<51>:I q<52>:I q<53>:I q<54>:I q<55>:I 
*.PININFO q<56>:I q<57>:I q<58>:I q<59>:I q<60>:I q<61>:I q<62>:I q<63>:I 
*.PININFO time<0>:I time<1>:I time<2>:I time<3>:I in1<0>:O in1<1>:O in1<2>:O 
*.PININFO in1<3>:O in1<4>:O in1<5>:O in1<6>:O in1<7>:O in1<8>:O in1<9>:O 
*.PININFO in1<10>:O in1<11>:O in1<12>:O in1<13>:O in1<14>:O in1<15>:O in2<0>:O 
*.PININFO in2<1>:O in2<2>:O in2<3>:O in2<4>:O in2<5>:O in2<6>:O in2<7>:O 
*.PININFO in2<8>:O in2<9>:O in2<10>:O in2<11>:O in2<12>:O in2<13>:O in2<14>:O 
*.PININFO in2<15>:O vdd:B vss:B
XI134 entime in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> 
+ in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> q<32> q<33> 
+ q<34> q<35> q<36> q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> 
+ q<46> q<47> q<48> q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> 
+ q<58> q<59> q<60> q<61> q<62> q<63> time<0> time<1> time<2> time<3> vdd vss 
+ / Tgenerate_array_8
XI133 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in2<0> 
+ in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> q<0> q<1> q<2> q<3> q<4> 
+ q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> q<15> q<16> q<17> 
+ q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> q<27> q<28> q<29> 
+ q<30> q<31> time<0> time<1> time<2> time<3> vdd vss / Tgenerate_array_8
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_32
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_32 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> 
+ in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> 
+ in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> 
+ in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in2<0> in2<1> in2<2> 
+ in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> 
+ in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> 
+ in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> 
+ in2<31> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> 
+ q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> 
+ q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> 
+ q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> 
+ q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> 
+ q<61> q<62> q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> 
+ q<73> q<74> q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> 
+ q<85> q<86> q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> 
+ q<97> q<98> q<99> q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> 
+ q<108> q<109> q<110> q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> 
+ q<119> q<120> q<121> q<122> q<123> q<124> q<125> q<126> q<127> time<0> 
+ time<1> time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO q<16>:I q<17>:I q<18>:I q<19>:I q<20>:I q<21>:I q<22>:I q<23>:I 
*.PININFO q<24>:I q<25>:I q<26>:I q<27>:I q<28>:I q<29>:I q<30>:I q<31>:I 
*.PININFO q<32>:I q<33>:I q<34>:I q<35>:I q<36>:I q<37>:I q<38>:I q<39>:I 
*.PININFO q<40>:I q<41>:I q<42>:I q<43>:I q<44>:I q<45>:I q<46>:I q<47>:I 
*.PININFO q<48>:I q<49>:I q<50>:I q<51>:I q<52>:I q<53>:I q<54>:I q<55>:I 
*.PININFO q<56>:I q<57>:I q<58>:I q<59>:I q<60>:I q<61>:I q<62>:I q<63>:I 
*.PININFO q<64>:I q<65>:I q<66>:I q<67>:I q<68>:I q<69>:I q<70>:I q<71>:I 
*.PININFO q<72>:I q<73>:I q<74>:I q<75>:I q<76>:I q<77>:I q<78>:I q<79>:I 
*.PININFO q<80>:I q<81>:I q<82>:I q<83>:I q<84>:I q<85>:I q<86>:I q<87>:I 
*.PININFO q<88>:I q<89>:I q<90>:I q<91>:I q<92>:I q<93>:I q<94>:I q<95>:I 
*.PININFO q<96>:I q<97>:I q<98>:I q<99>:I q<100>:I q<101>:I q<102>:I q<103>:I 
*.PININFO q<104>:I q<105>:I q<106>:I q<107>:I q<108>:I q<109>:I q<110>:I 
*.PININFO q<111>:I q<112>:I q<113>:I q<114>:I q<115>:I q<116>:I q<117>:I 
*.PININFO q<118>:I q<119>:I q<120>:I q<121>:I q<122>:I q<123>:I q<124>:I 
*.PININFO q<125>:I q<126>:I q<127>:I time<0>:I time<1>:I time<2>:I time<3>:I 
*.PININFO in1<0>:O in1<1>:O in1<2>:O in1<3>:O in1<4>:O in1<5>:O in1<6>:O 
*.PININFO in1<7>:O in1<8>:O in1<9>:O in1<10>:O in1<11>:O in1<12>:O in1<13>:O 
*.PININFO in1<14>:O in1<15>:O in1<16>:O in1<17>:O in1<18>:O in1<19>:O 
*.PININFO in1<20>:O in1<21>:O in1<22>:O in1<23>:O in1<24>:O in1<25>:O 
*.PININFO in1<26>:O in1<27>:O in1<28>:O in1<29>:O in1<30>:O in1<31>:O in2<0>:O 
*.PININFO in2<1>:O in2<2>:O in2<3>:O in2<4>:O in2<5>:O in2<6>:O in2<7>:O 
*.PININFO in2<8>:O in2<9>:O in2<10>:O in2<11>:O in2<12>:O in2<13>:O in2<14>:O 
*.PININFO in2<15>:O in2<16>:O in2<17>:O in2<18>:O in2<19>:O in2<20>:O 
*.PININFO in2<21>:O in2<22>:O in2<23>:O in2<24>:O in2<25>:O in2<26>:O 
*.PININFO in2<27>:O in2<28>:O in2<29>:O in2<30>:O in2<31>:O vdd:B vss:B
XI135 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> 
+ in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in2<0> in2<1> in2<2> 
+ in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> 
+ in2<13> in2<14> in2<15> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> 
+ q<10> q<11> q<12> q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> 
+ q<22> q<23> q<24> q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> 
+ q<34> q<35> q<36> q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> 
+ q<46> q<47> q<48> q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> 
+ q<58> q<59> q<60> q<61> q<62> q<63> time<0> time<1> time<2> time<3> vdd vss 
+ / Tgenerate_array_16
XI136 entime in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> 
+ in1<24> in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in2<16> 
+ in2<17> in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> 
+ in2<26> in2<27> in2<28> in2<29> in2<30> in2<31> q<64> q<65> q<66> q<67> 
+ q<68> q<69> q<70> q<71> q<72> q<73> q<74> q<75> q<76> q<77> q<78> q<79> 
+ q<80> q<81> q<82> q<83> q<84> q<85> q<86> q<87> q<88> q<89> q<90> q<91> 
+ q<92> q<93> q<94> q<95> q<96> q<97> q<98> q<99> q<100> q<101> q<102> q<103> 
+ q<104> q<105> q<106> q<107> q<108> q<109> q<110> q<111> q<112> q<113> q<114> 
+ q<115> q<116> q<117> q<118> q<119> q<120> q<121> q<122> q<123> q<124> q<125> 
+ q<126> q<127> time<0> time<1> time<2> time<3> vdd vss / Tgenerate_array_16
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_64
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_64 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> 
+ in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> 
+ in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> 
+ in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> 
+ in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> 
+ in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> 
+ in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> 
+ in1<61> in1<62> in1<63> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> 
+ in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> 
+ in2<17> in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> 
+ in2<26> in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> 
+ in2<35> in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> 
+ in2<44> in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> 
+ in2<53> in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> 
+ in2<62> in2<63> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> 
+ q<11> q<12> q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> 
+ q<23> q<24> q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> 
+ q<35> q<36> q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> 
+ q<47> q<48> q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> 
+ q<59> q<60> q<61> q<62> q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> 
+ q<71> q<72> q<73> q<74> q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> 
+ q<83> q<84> q<85> q<86> q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> 
+ q<95> q<96> q<97> q<98> q<99> q<100> q<101> q<102> q<103> q<104> q<105> 
+ q<106> q<107> q<108> q<109> q<110> q<111> q<112> q<113> q<114> q<115> q<116> 
+ q<117> q<118> q<119> q<120> q<121> q<122> q<123> q<124> q<125> q<126> q<127> 
+ q<128> q<129> q<130> q<131> q<132> q<133> q<134> q<135> q<136> q<137> q<138> 
+ q<139> q<140> q<141> q<142> q<143> q<144> q<145> q<146> q<147> q<148> q<149> 
+ q<150> q<151> q<152> q<153> q<154> q<155> q<156> q<157> q<158> q<159> q<160> 
+ q<161> q<162> q<163> q<164> q<165> q<166> q<167> q<168> q<169> q<170> q<171> 
+ q<172> q<173> q<174> q<175> q<176> q<177> q<178> q<179> q<180> q<181> q<182> 
+ q<183> q<184> q<185> q<186> q<187> q<188> q<189> q<190> q<191> q<192> q<193> 
+ q<194> q<195> q<196> q<197> q<198> q<199> q<200> q<201> q<202> q<203> q<204> 
+ q<205> q<206> q<207> q<208> q<209> q<210> q<211> q<212> q<213> q<214> q<215> 
+ q<216> q<217> q<218> q<219> q<220> q<221> q<222> q<223> q<224> q<225> q<226> 
+ q<227> q<228> q<229> q<230> q<231> q<232> q<233> q<234> q<235> q<236> q<237> 
+ q<238> q<239> q<240> q<241> q<242> q<243> q<244> q<245> q<246> q<247> q<248> 
+ q<249> q<250> q<251> q<252> q<253> q<254> q<255> time<0> time<1> time<2> 
+ time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO q<16>:I q<17>:I q<18>:I q<19>:I q<20>:I q<21>:I q<22>:I q<23>:I 
*.PININFO q<24>:I q<25>:I q<26>:I q<27>:I q<28>:I q<29>:I q<30>:I q<31>:I 
*.PININFO q<32>:I q<33>:I q<34>:I q<35>:I q<36>:I q<37>:I q<38>:I q<39>:I 
*.PININFO q<40>:I q<41>:I q<42>:I q<43>:I q<44>:I q<45>:I q<46>:I q<47>:I 
*.PININFO q<48>:I q<49>:I q<50>:I q<51>:I q<52>:I q<53>:I q<54>:I q<55>:I 
*.PININFO q<56>:I q<57>:I q<58>:I q<59>:I q<60>:I q<61>:I q<62>:I q<63>:I 
*.PININFO q<64>:I q<65>:I q<66>:I q<67>:I q<68>:I q<69>:I q<70>:I q<71>:I 
*.PININFO q<72>:I q<73>:I q<74>:I q<75>:I q<76>:I q<77>:I q<78>:I q<79>:I 
*.PININFO q<80>:I q<81>:I q<82>:I q<83>:I q<84>:I q<85>:I q<86>:I q<87>:I 
*.PININFO q<88>:I q<89>:I q<90>:I q<91>:I q<92>:I q<93>:I q<94>:I q<95>:I 
*.PININFO q<96>:I q<97>:I q<98>:I q<99>:I q<100>:I q<101>:I q<102>:I q<103>:I 
*.PININFO q<104>:I q<105>:I q<106>:I q<107>:I q<108>:I q<109>:I q<110>:I 
*.PININFO q<111>:I q<112>:I q<113>:I q<114>:I q<115>:I q<116>:I q<117>:I 
*.PININFO q<118>:I q<119>:I q<120>:I q<121>:I q<122>:I q<123>:I q<124>:I 
*.PININFO q<125>:I q<126>:I q<127>:I q<128>:I q<129>:I q<130>:I q<131>:I 
*.PININFO q<132>:I q<133>:I q<134>:I q<135>:I q<136>:I q<137>:I q<138>:I 
*.PININFO q<139>:I q<140>:I q<141>:I q<142>:I q<143>:I q<144>:I q<145>:I 
*.PININFO q<146>:I q<147>:I q<148>:I q<149>:I q<150>:I q<151>:I q<152>:I 
*.PININFO q<153>:I q<154>:I q<155>:I q<156>:I q<157>:I q<158>:I q<159>:I 
*.PININFO q<160>:I q<161>:I q<162>:I q<163>:I q<164>:I q<165>:I q<166>:I 
*.PININFO q<167>:I q<168>:I q<169>:I q<170>:I q<171>:I q<172>:I q<173>:I 
*.PININFO q<174>:I q<175>:I q<176>:I q<177>:I q<178>:I q<179>:I q<180>:I 
*.PININFO q<181>:I q<182>:I q<183>:I q<184>:I q<185>:I q<186>:I q<187>:I 
*.PININFO q<188>:I q<189>:I q<190>:I q<191>:I q<192>:I q<193>:I q<194>:I 
*.PININFO q<195>:I q<196>:I q<197>:I q<198>:I q<199>:I q<200>:I q<201>:I 
*.PININFO q<202>:I q<203>:I q<204>:I q<205>:I q<206>:I q<207>:I q<208>:I 
*.PININFO q<209>:I q<210>:I q<211>:I q<212>:I q<213>:I q<214>:I q<215>:I 
*.PININFO q<216>:I q<217>:I q<218>:I q<219>:I q<220>:I q<221>:I q<222>:I 
*.PININFO q<223>:I q<224>:I q<225>:I q<226>:I q<227>:I q<228>:I q<229>:I 
*.PININFO q<230>:I q<231>:I q<232>:I q<233>:I q<234>:I q<235>:I q<236>:I 
*.PININFO q<237>:I q<238>:I q<239>:I q<240>:I q<241>:I q<242>:I q<243>:I 
*.PININFO q<244>:I q<245>:I q<246>:I q<247>:I q<248>:I q<249>:I q<250>:I 
*.PININFO q<251>:I q<252>:I q<253>:I q<254>:I q<255>:I time<0>:I time<1>:I 
*.PININFO time<2>:I time<3>:I in1<0>:O in1<1>:O in1<2>:O in1<3>:O in1<4>:O 
*.PININFO in1<5>:O in1<6>:O in1<7>:O in1<8>:O in1<9>:O in1<10>:O in1<11>:O 
*.PININFO in1<12>:O in1<13>:O in1<14>:O in1<15>:O in1<16>:O in1<17>:O 
*.PININFO in1<18>:O in1<19>:O in1<20>:O in1<21>:O in1<22>:O in1<23>:O 
*.PININFO in1<24>:O in1<25>:O in1<26>:O in1<27>:O in1<28>:O in1<29>:O 
*.PININFO in1<30>:O in1<31>:O in1<32>:O in1<33>:O in1<34>:O in1<35>:O 
*.PININFO in1<36>:O in1<37>:O in1<38>:O in1<39>:O in1<40>:O in1<41>:O 
*.PININFO in1<42>:O in1<43>:O in1<44>:O in1<45>:O in1<46>:O in1<47>:O 
*.PININFO in1<48>:O in1<49>:O in1<50>:O in1<51>:O in1<52>:O in1<53>:O 
*.PININFO in1<54>:O in1<55>:O in1<56>:O in1<57>:O in1<58>:O in1<59>:O 
*.PININFO in1<60>:O in1<61>:O in1<62>:O in1<63>:O in2<0>:O in2<1>:O in2<2>:O 
*.PININFO in2<3>:O in2<4>:O in2<5>:O in2<6>:O in2<7>:O in2<8>:O in2<9>:O 
*.PININFO in2<10>:O in2<11>:O in2<12>:O in2<13>:O in2<14>:O in2<15>:O 
*.PININFO in2<16>:O in2<17>:O in2<18>:O in2<19>:O in2<20>:O in2<21>:O 
*.PININFO in2<22>:O in2<23>:O in2<24>:O in2<25>:O in2<26>:O in2<27>:O 
*.PININFO in2<28>:O in2<29>:O in2<30>:O in2<31>:O in2<32>:O in2<33>:O 
*.PININFO in2<34>:O in2<35>:O in2<36>:O in2<37>:O in2<38>:O in2<39>:O 
*.PININFO in2<40>:O in2<41>:O in2<42>:O in2<43>:O in2<44>:O in2<45>:O 
*.PININFO in2<46>:O in2<47>:O in2<48>:O in2<49>:O in2<50>:O in2<51>:O 
*.PININFO in2<52>:O in2<53>:O in2<54>:O in2<55>:O in2<56>:O in2<57>:O 
*.PININFO in2<58>:O in2<59>:O in2<60>:O in2<61>:O in2<62>:O in2<63>:O vdd:B 
*.PININFO vss:B
XI25<0> time<0> net013<0> vdd vss / inv4
XI25<1> time<1> net013<1> vdd vss / inv4
XI25<2> time<2> net013<2> vdd vss / inv4
XI25<3> time<3> net013<3> vdd vss / inv4
XI3 entime net011 vdd vss / inv4
XI138 entimeb in1<32> in1<33> in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> 
+ in1<40> in1<41> in1<42> in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> 
+ in1<49> in1<50> in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> 
+ in1<58> in1<59> in1<60> in1<61> in1<62> in1<63> in2<32> in2<33> in2<34> 
+ in2<35> in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> 
+ in2<44> in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> 
+ in2<53> in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> 
+ in2<62> in2<63> q<128> q<129> q<130> q<131> q<132> q<133> q<134> q<135> 
+ q<136> q<137> q<138> q<139> q<140> q<141> q<142> q<143> q<144> q<145> q<146> 
+ q<147> q<148> q<149> q<150> q<151> q<152> q<153> q<154> q<155> q<156> q<157> 
+ q<158> q<159> q<160> q<161> q<162> q<163> q<164> q<165> q<166> q<167> q<168> 
+ q<169> q<170> q<171> q<172> q<173> q<174> q<175> q<176> q<177> q<178> q<179> 
+ q<180> q<181> q<182> q<183> q<184> q<185> q<186> q<187> q<188> q<189> q<190> 
+ q<191> q<192> q<193> q<194> q<195> q<196> q<197> q<198> q<199> q<200> q<201> 
+ q<202> q<203> q<204> q<205> q<206> q<207> q<208> q<209> q<210> q<211> q<212> 
+ q<213> q<214> q<215> q<216> q<217> q<218> q<219> q<220> q<221> q<222> q<223> 
+ q<224> q<225> q<226> q<227> q<228> q<229> q<230> q<231> q<232> q<233> q<234> 
+ q<235> q<236> q<237> q<238> q<239> q<240> q<241> q<242> q<243> q<244> q<245> 
+ q<246> q<247> q<248> q<249> q<250> q<251> q<252> q<253> q<254> q<255> 
+ timeb<0> timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate_array_32
XI137 entimeb in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> 
+ in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> in1<17> 
+ in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> in1<26> 
+ in1<27> in1<28> in1<29> in1<30> in1<31> in2<0> in2<1> in2<2> in2<3> in2<4> 
+ in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> 
+ in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> 
+ in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> in2<31> q<0> q<1> 
+ q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> q<15> 
+ q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> q<27> 
+ q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> q<37> q<38> q<39> 
+ q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> q<49> q<50> q<51> 
+ q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> q<61> q<62> q<63> 
+ q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> q<73> q<74> q<75> 
+ q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> q<85> q<86> q<87> 
+ q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> q<97> q<98> q<99> 
+ q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> q<108> q<109> q<110> 
+ q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> q<119> q<120> q<121> 
+ q<122> q<123> q<124> q<125> q<126> q<127> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate_array_32
XI2 net011 entimeb vdd vss / inv8
XI1<0> net013<0> timeb<0> vdd vss / inv8
XI1<1> net013<1> timeb<1> vdd vss / inv8
XI1<2> net013<2> timeb<2> vdd vss / inv8
XI1<3> net013<3> timeb<3> vdd vss / inv8
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate_array_128
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate_array_128 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> 
+ in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> 
+ in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> 
+ in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> 
+ in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> 
+ in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> 
+ in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> 
+ in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> 
+ in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> 
+ in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> 
+ in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> 
+ in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> 
+ in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> 
+ in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> 
+ in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> 
+ in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> 
+ in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> 
+ in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> 
+ in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> 
+ in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> 
+ in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> 
+ in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> 
+ in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> 
+ in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> 
+ in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> 
+ in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> 
+ in2<102> in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> 
+ in2<110> in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> 
+ in2<118> in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> 
+ in2<126> in2<127> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> 
+ q<11> q<12> q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> 
+ q<23> q<24> q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> 
+ q<35> q<36> q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> 
+ q<47> q<48> q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> 
+ q<59> q<60> q<61> q<62> q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> 
+ q<71> q<72> q<73> q<74> q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> 
+ q<83> q<84> q<85> q<86> q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> 
+ q<95> q<96> q<97> q<98> q<99> q<100> q<101> q<102> q<103> q<104> q<105> 
+ q<106> q<107> q<108> q<109> q<110> q<111> q<112> q<113> q<114> q<115> q<116> 
+ q<117> q<118> q<119> q<120> q<121> q<122> q<123> q<124> q<125> q<126> q<127> 
+ q<128> q<129> q<130> q<131> q<132> q<133> q<134> q<135> q<136> q<137> q<138> 
+ q<139> q<140> q<141> q<142> q<143> q<144> q<145> q<146> q<147> q<148> q<149> 
+ q<150> q<151> q<152> q<153> q<154> q<155> q<156> q<157> q<158> q<159> q<160> 
+ q<161> q<162> q<163> q<164> q<165> q<166> q<167> q<168> q<169> q<170> q<171> 
+ q<172> q<173> q<174> q<175> q<176> q<177> q<178> q<179> q<180> q<181> q<182> 
+ q<183> q<184> q<185> q<186> q<187> q<188> q<189> q<190> q<191> q<192> q<193> 
+ q<194> q<195> q<196> q<197> q<198> q<199> q<200> q<201> q<202> q<203> q<204> 
+ q<205> q<206> q<207> q<208> q<209> q<210> q<211> q<212> q<213> q<214> q<215> 
+ q<216> q<217> q<218> q<219> q<220> q<221> q<222> q<223> q<224> q<225> q<226> 
+ q<227> q<228> q<229> q<230> q<231> q<232> q<233> q<234> q<235> q<236> q<237> 
+ q<238> q<239> q<240> q<241> q<242> q<243> q<244> q<245> q<246> q<247> q<248> 
+ q<249> q<250> q<251> q<252> q<253> q<254> q<255> q<256> q<257> q<258> q<259> 
+ q<260> q<261> q<262> q<263> q<264> q<265> q<266> q<267> q<268> q<269> q<270> 
+ q<271> q<272> q<273> q<274> q<275> q<276> q<277> q<278> q<279> q<280> q<281> 
+ q<282> q<283> q<284> q<285> q<286> q<287> q<288> q<289> q<290> q<291> q<292> 
+ q<293> q<294> q<295> q<296> q<297> q<298> q<299> q<300> q<301> q<302> q<303> 
+ q<304> q<305> q<306> q<307> q<308> q<309> q<310> q<311> q<312> q<313> q<314> 
+ q<315> q<316> q<317> q<318> q<319> q<320> q<321> q<322> q<323> q<324> q<325> 
+ q<326> q<327> q<328> q<329> q<330> q<331> q<332> q<333> q<334> q<335> q<336> 
+ q<337> q<338> q<339> q<340> q<341> q<342> q<343> q<344> q<345> q<346> q<347> 
+ q<348> q<349> q<350> q<351> q<352> q<353> q<354> q<355> q<356> q<357> q<358> 
+ q<359> q<360> q<361> q<362> q<363> q<364> q<365> q<366> q<367> q<368> q<369> 
+ q<370> q<371> q<372> q<373> q<374> q<375> q<376> q<377> q<378> q<379> q<380> 
+ q<381> q<382> q<383> q<384> q<385> q<386> q<387> q<388> q<389> q<390> q<391> 
+ q<392> q<393> q<394> q<395> q<396> q<397> q<398> q<399> q<400> q<401> q<402> 
+ q<403> q<404> q<405> q<406> q<407> q<408> q<409> q<410> q<411> q<412> q<413> 
+ q<414> q<415> q<416> q<417> q<418> q<419> q<420> q<421> q<422> q<423> q<424> 
+ q<425> q<426> q<427> q<428> q<429> q<430> q<431> q<432> q<433> q<434> q<435> 
+ q<436> q<437> q<438> q<439> q<440> q<441> q<442> q<443> q<444> q<445> q<446> 
+ q<447> q<448> q<449> q<450> q<451> q<452> q<453> q<454> q<455> q<456> q<457> 
+ q<458> q<459> q<460> q<461> q<462> q<463> q<464> q<465> q<466> q<467> q<468> 
+ q<469> q<470> q<471> q<472> q<473> q<474> q<475> q<476> q<477> q<478> q<479> 
+ q<480> q<481> q<482> q<483> q<484> q<485> q<486> q<487> q<488> q<489> q<490> 
+ q<491> q<492> q<493> q<494> q<495> q<496> q<497> q<498> q<499> q<500> q<501> 
+ q<502> q<503> q<504> q<505> q<506> q<507> q<508> q<509> q<510> q<511> 
+ time<0> time<1> time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO q<16>:I q<17>:I q<18>:I q<19>:I q<20>:I q<21>:I q<22>:I q<23>:I 
*.PININFO q<24>:I q<25>:I q<26>:I q<27>:I q<28>:I q<29>:I q<30>:I q<31>:I 
*.PININFO q<32>:I q<33>:I q<34>:I q<35>:I q<36>:I q<37>:I q<38>:I q<39>:I 
*.PININFO q<40>:I q<41>:I q<42>:I q<43>:I q<44>:I q<45>:I q<46>:I q<47>:I 
*.PININFO q<48>:I q<49>:I q<50>:I q<51>:I q<52>:I q<53>:I q<54>:I q<55>:I 
*.PININFO q<56>:I q<57>:I q<58>:I q<59>:I q<60>:I q<61>:I q<62>:I q<63>:I 
*.PININFO q<64>:I q<65>:I q<66>:I q<67>:I q<68>:I q<69>:I q<70>:I q<71>:I 
*.PININFO q<72>:I q<73>:I q<74>:I q<75>:I q<76>:I q<77>:I q<78>:I q<79>:I 
*.PININFO q<80>:I q<81>:I q<82>:I q<83>:I q<84>:I q<85>:I q<86>:I q<87>:I 
*.PININFO q<88>:I q<89>:I q<90>:I q<91>:I q<92>:I q<93>:I q<94>:I q<95>:I 
*.PININFO q<96>:I q<97>:I q<98>:I q<99>:I q<100>:I q<101>:I q<102>:I q<103>:I 
*.PININFO q<104>:I q<105>:I q<106>:I q<107>:I q<108>:I q<109>:I q<110>:I 
*.PININFO q<111>:I q<112>:I q<113>:I q<114>:I q<115>:I q<116>:I q<117>:I 
*.PININFO q<118>:I q<119>:I q<120>:I q<121>:I q<122>:I q<123>:I q<124>:I 
*.PININFO q<125>:I q<126>:I q<127>:I q<128>:I q<129>:I q<130>:I q<131>:I 
*.PININFO q<132>:I q<133>:I q<134>:I q<135>:I q<136>:I q<137>:I q<138>:I 
*.PININFO q<139>:I q<140>:I q<141>:I q<142>:I q<143>:I q<144>:I q<145>:I 
*.PININFO q<146>:I q<147>:I q<148>:I q<149>:I q<150>:I q<151>:I q<152>:I 
*.PININFO q<153>:I q<154>:I q<155>:I q<156>:I q<157>:I q<158>:I q<159>:I 
*.PININFO q<160>:I q<161>:I q<162>:I q<163>:I q<164>:I q<165>:I q<166>:I 
*.PININFO q<167>:I q<168>:I q<169>:I q<170>:I q<171>:I q<172>:I q<173>:I 
*.PININFO q<174>:I q<175>:I q<176>:I q<177>:I q<178>:I q<179>:I q<180>:I 
*.PININFO q<181>:I q<182>:I q<183>:I q<184>:I q<185>:I q<186>:I q<187>:I 
*.PININFO q<188>:I q<189>:I q<190>:I q<191>:I q<192>:I q<193>:I q<194>:I 
*.PININFO q<195>:I q<196>:I q<197>:I q<198>:I q<199>:I q<200>:I q<201>:I 
*.PININFO q<202>:I q<203>:I q<204>:I q<205>:I q<206>:I q<207>:I q<208>:I 
*.PININFO q<209>:I q<210>:I q<211>:I q<212>:I q<213>:I q<214>:I q<215>:I 
*.PININFO q<216>:I q<217>:I q<218>:I q<219>:I q<220>:I q<221>:I q<222>:I 
*.PININFO q<223>:I q<224>:I q<225>:I q<226>:I q<227>:I q<228>:I q<229>:I 
*.PININFO q<230>:I q<231>:I q<232>:I q<233>:I q<234>:I q<235>:I q<236>:I 
*.PININFO q<237>:I q<238>:I q<239>:I q<240>:I q<241>:I q<242>:I q<243>:I 
*.PININFO q<244>:I q<245>:I q<246>:I q<247>:I q<248>:I q<249>:I q<250>:I 
*.PININFO q<251>:I q<252>:I q<253>:I q<254>:I q<255>:I q<256>:I q<257>:I 
*.PININFO q<258>:I q<259>:I q<260>:I q<261>:I q<262>:I q<263>:I q<264>:I 
*.PININFO q<265>:I q<266>:I q<267>:I q<268>:I q<269>:I q<270>:I q<271>:I 
*.PININFO q<272>:I q<273>:I q<274>:I q<275>:I q<276>:I q<277>:I q<278>:I 
*.PININFO q<279>:I q<280>:I q<281>:I q<282>:I q<283>:I q<284>:I q<285>:I 
*.PININFO q<286>:I q<287>:I q<288>:I q<289>:I q<290>:I q<291>:I q<292>:I 
*.PININFO q<293>:I q<294>:I q<295>:I q<296>:I q<297>:I q<298>:I q<299>:I 
*.PININFO q<300>:I q<301>:I q<302>:I q<303>:I q<304>:I q<305>:I q<306>:I 
*.PININFO q<307>:I q<308>:I q<309>:I q<310>:I q<311>:I q<312>:I q<313>:I 
*.PININFO q<314>:I q<315>:I q<316>:I q<317>:I q<318>:I q<319>:I q<320>:I 
*.PININFO q<321>:I q<322>:I q<323>:I q<324>:I q<325>:I q<326>:I q<327>:I 
*.PININFO q<328>:I q<329>:I q<330>:I q<331>:I q<332>:I q<333>:I q<334>:I 
*.PININFO q<335>:I q<336>:I q<337>:I q<338>:I q<339>:I q<340>:I q<341>:I 
*.PININFO q<342>:I q<343>:I q<344>:I q<345>:I q<346>:I q<347>:I q<348>:I 
*.PININFO q<349>:I q<350>:I q<351>:I q<352>:I q<353>:I q<354>:I q<355>:I 
*.PININFO q<356>:I q<357>:I q<358>:I q<359>:I q<360>:I q<361>:I q<362>:I 
*.PININFO q<363>:I q<364>:I q<365>:I q<366>:I q<367>:I q<368>:I q<369>:I 
*.PININFO q<370>:I q<371>:I q<372>:I q<373>:I q<374>:I q<375>:I q<376>:I 
*.PININFO q<377>:I q<378>:I q<379>:I q<380>:I q<381>:I q<382>:I q<383>:I 
*.PININFO q<384>:I q<385>:I q<386>:I q<387>:I q<388>:I q<389>:I q<390>:I 
*.PININFO q<391>:I q<392>:I q<393>:I q<394>:I q<395>:I q<396>:I q<397>:I 
*.PININFO q<398>:I q<399>:I q<400>:I q<401>:I q<402>:I q<403>:I q<404>:I 
*.PININFO q<405>:I q<406>:I q<407>:I q<408>:I q<409>:I q<410>:I q<411>:I 
*.PININFO q<412>:I q<413>:I q<414>:I q<415>:I q<416>:I q<417>:I q<418>:I 
*.PININFO q<419>:I q<420>:I q<421>:I q<422>:I q<423>:I q<424>:I q<425>:I 
*.PININFO q<426>:I q<427>:I q<428>:I q<429>:I q<430>:I q<431>:I q<432>:I 
*.PININFO q<433>:I q<434>:I q<435>:I q<436>:I q<437>:I q<438>:I q<439>:I 
*.PININFO q<440>:I q<441>:I q<442>:I q<443>:I q<444>:I q<445>:I q<446>:I 
*.PININFO q<447>:I q<448>:I q<449>:I q<450>:I q<451>:I q<452>:I q<453>:I 
*.PININFO q<454>:I q<455>:I q<456>:I q<457>:I q<458>:I q<459>:I q<460>:I 
*.PININFO q<461>:I q<462>:I q<463>:I q<464>:I q<465>:I q<466>:I q<467>:I 
*.PININFO q<468>:I q<469>:I q<470>:I q<471>:I q<472>:I q<473>:I q<474>:I 
*.PININFO q<475>:I q<476>:I q<477>:I q<478>:I q<479>:I q<480>:I q<481>:I 
*.PININFO q<482>:I q<483>:I q<484>:I q<485>:I q<486>:I q<487>:I q<488>:I 
*.PININFO q<489>:I q<490>:I q<491>:I q<492>:I q<493>:I q<494>:I q<495>:I 
*.PININFO q<496>:I q<497>:I q<498>:I q<499>:I q<500>:I q<501>:I q<502>:I 
*.PININFO q<503>:I q<504>:I q<505>:I q<506>:I q<507>:I q<508>:I q<509>:I 
*.PININFO q<510>:I q<511>:I time<0>:I time<1>:I time<2>:I time<3>:I in1<0>:O 
*.PININFO in1<1>:O in1<2>:O in1<3>:O in1<4>:O in1<5>:O in1<6>:O in1<7>:O 
*.PININFO in1<8>:O in1<9>:O in1<10>:O in1<11>:O in1<12>:O in1<13>:O in1<14>:O 
*.PININFO in1<15>:O in1<16>:O in1<17>:O in1<18>:O in1<19>:O in1<20>:O 
*.PININFO in1<21>:O in1<22>:O in1<23>:O in1<24>:O in1<25>:O in1<26>:O 
*.PININFO in1<27>:O in1<28>:O in1<29>:O in1<30>:O in1<31>:O in1<32>:O 
*.PININFO in1<33>:O in1<34>:O in1<35>:O in1<36>:O in1<37>:O in1<38>:O 
*.PININFO in1<39>:O in1<40>:O in1<41>:O in1<42>:O in1<43>:O in1<44>:O 
*.PININFO in1<45>:O in1<46>:O in1<47>:O in1<48>:O in1<49>:O in1<50>:O 
*.PININFO in1<51>:O in1<52>:O in1<53>:O in1<54>:O in1<55>:O in1<56>:O 
*.PININFO in1<57>:O in1<58>:O in1<59>:O in1<60>:O in1<61>:O in1<62>:O 
*.PININFO in1<63>:O in1<64>:O in1<65>:O in1<66>:O in1<67>:O in1<68>:O 
*.PININFO in1<69>:O in1<70>:O in1<71>:O in1<72>:O in1<73>:O in1<74>:O 
*.PININFO in1<75>:O in1<76>:O in1<77>:O in1<78>:O in1<79>:O in1<80>:O 
*.PININFO in1<81>:O in1<82>:O in1<83>:O in1<84>:O in1<85>:O in1<86>:O 
*.PININFO in1<87>:O in1<88>:O in1<89>:O in1<90>:O in1<91>:O in1<92>:O 
*.PININFO in1<93>:O in1<94>:O in1<95>:O in1<96>:O in1<97>:O in1<98>:O 
*.PININFO in1<99>:O in1<100>:O in1<101>:O in1<102>:O in1<103>:O in1<104>:O 
*.PININFO in1<105>:O in1<106>:O in1<107>:O in1<108>:O in1<109>:O in1<110>:O 
*.PININFO in1<111>:O in1<112>:O in1<113>:O in1<114>:O in1<115>:O in1<116>:O 
*.PININFO in1<117>:O in1<118>:O in1<119>:O in1<120>:O in1<121>:O in1<122>:O 
*.PININFO in1<123>:O in1<124>:O in1<125>:O in1<126>:O in1<127>:O in2<0>:O 
*.PININFO in2<1>:O in2<2>:O in2<3>:O in2<4>:O in2<5>:O in2<6>:O in2<7>:O 
*.PININFO in2<8>:O in2<9>:O in2<10>:O in2<11>:O in2<12>:O in2<13>:O in2<14>:O 
*.PININFO in2<15>:O in2<16>:O in2<17>:O in2<18>:O in2<19>:O in2<20>:O 
*.PININFO in2<21>:O in2<22>:O in2<23>:O in2<24>:O in2<25>:O in2<26>:O 
*.PININFO in2<27>:O in2<28>:O in2<29>:O in2<30>:O in2<31>:O in2<32>:O 
*.PININFO in2<33>:O in2<34>:O in2<35>:O in2<36>:O in2<37>:O in2<38>:O 
*.PININFO in2<39>:O in2<40>:O in2<41>:O in2<42>:O in2<43>:O in2<44>:O 
*.PININFO in2<45>:O in2<46>:O in2<47>:O in2<48>:O in2<49>:O in2<50>:O 
*.PININFO in2<51>:O in2<52>:O in2<53>:O in2<54>:O in2<55>:O in2<56>:O 
*.PININFO in2<57>:O in2<58>:O in2<59>:O in2<60>:O in2<61>:O in2<62>:O 
*.PININFO in2<63>:O in2<64>:O in2<65>:O in2<66>:O in2<67>:O in2<68>:O 
*.PININFO in2<69>:O in2<70>:O in2<71>:O in2<72>:O in2<73>:O in2<74>:O 
*.PININFO in2<75>:O in2<76>:O in2<77>:O in2<78>:O in2<79>:O in2<80>:O 
*.PININFO in2<81>:O in2<82>:O in2<83>:O in2<84>:O in2<85>:O in2<86>:O 
*.PININFO in2<87>:O in2<88>:O in2<89>:O in2<90>:O in2<91>:O in2<92>:O 
*.PININFO in2<93>:O in2<94>:O in2<95>:O in2<96>:O in2<97>:O in2<98>:O 
*.PININFO in2<99>:O in2<100>:O in2<101>:O in2<102>:O in2<103>:O in2<104>:O 
*.PININFO in2<105>:O in2<106>:O in2<107>:O in2<108>:O in2<109>:O in2<110>:O 
*.PININFO in2<111>:O in2<112>:O in2<113>:O in2<114>:O in2<115>:O in2<116>:O 
*.PININFO in2<117>:O in2<118>:O in2<119>:O in2<120>:O in2<121>:O in2<122>:O 
*.PININFO in2<123>:O in2<124>:O in2<125>:O in2<126>:O in2<127>:O vdd:B vss:B
XI130 entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> 
+ in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> in1<17> 
+ in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> in1<26> 
+ in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> in1<35> 
+ in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> in1<44> 
+ in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> in1<53> 
+ in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> in1<62> 
+ in1<63> in2<0> in2<1> in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> 
+ in2<9> in2<10> in2<11> in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> 
+ in2<18> in2<19> in2<20> in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> 
+ in2<27> in2<28> in2<29> in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> 
+ in2<36> in2<37> in2<38> in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> 
+ in2<45> in2<46> in2<47> in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> 
+ in2<54> in2<55> in2<56> in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> 
+ in2<63> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> 
+ q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> 
+ q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> 
+ q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> 
+ q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> 
+ q<61> q<62> q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> 
+ q<73> q<74> q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> 
+ q<85> q<86> q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> 
+ q<97> q<98> q<99> q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> 
+ q<108> q<109> q<110> q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> 
+ q<119> q<120> q<121> q<122> q<123> q<124> q<125> q<126> q<127> q<128> q<129> 
+ q<130> q<131> q<132> q<133> q<134> q<135> q<136> q<137> q<138> q<139> q<140> 
+ q<141> q<142> q<143> q<144> q<145> q<146> q<147> q<148> q<149> q<150> q<151> 
+ q<152> q<153> q<154> q<155> q<156> q<157> q<158> q<159> q<160> q<161> q<162> 
+ q<163> q<164> q<165> q<166> q<167> q<168> q<169> q<170> q<171> q<172> q<173> 
+ q<174> q<175> q<176> q<177> q<178> q<179> q<180> q<181> q<182> q<183> q<184> 
+ q<185> q<186> q<187> q<188> q<189> q<190> q<191> q<192> q<193> q<194> q<195> 
+ q<196> q<197> q<198> q<199> q<200> q<201> q<202> q<203> q<204> q<205> q<206> 
+ q<207> q<208> q<209> q<210> q<211> q<212> q<213> q<214> q<215> q<216> q<217> 
+ q<218> q<219> q<220> q<221> q<222> q<223> q<224> q<225> q<226> q<227> q<228> 
+ q<229> q<230> q<231> q<232> q<233> q<234> q<235> q<236> q<237> q<238> q<239> 
+ q<240> q<241> q<242> q<243> q<244> q<245> q<246> q<247> q<248> q<249> q<250> 
+ q<251> q<252> q<253> q<254> q<255> time<0> time<1> time<2> time<3> vdd vss / 
+ Tgenerate_array_64
XI131 entime in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> in1<71> 
+ in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> in1<80> 
+ in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> in1<89> 
+ in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> in1<98> 
+ in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> in1<106> 
+ in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> in1<113> in1<114> 
+ in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> in1<122> 
+ in1<123> in1<124> in1<125> in1<126> in1<127> in2<64> in2<65> in2<66> in2<67> 
+ in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> in2<76> 
+ in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> in2<84> in2<85> 
+ in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> in2<94> 
+ in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> in2<102> in2<103> 
+ in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> in2<110> in2<111> 
+ in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> in2<118> in2<119> 
+ in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> in2<126> in2<127> 
+ q<256> q<257> q<258> q<259> q<260> q<261> q<262> q<263> q<264> q<265> q<266> 
+ q<267> q<268> q<269> q<270> q<271> q<272> q<273> q<274> q<275> q<276> q<277> 
+ q<278> q<279> q<280> q<281> q<282> q<283> q<284> q<285> q<286> q<287> q<288> 
+ q<289> q<290> q<291> q<292> q<293> q<294> q<295> q<296> q<297> q<298> q<299> 
+ q<300> q<301> q<302> q<303> q<304> q<305> q<306> q<307> q<308> q<309> q<310> 
+ q<311> q<312> q<313> q<314> q<315> q<316> q<317> q<318> q<319> q<320> q<321> 
+ q<322> q<323> q<324> q<325> q<326> q<327> q<328> q<329> q<330> q<331> q<332> 
+ q<333> q<334> q<335> q<336> q<337> q<338> q<339> q<340> q<341> q<342> q<343> 
+ q<344> q<345> q<346> q<347> q<348> q<349> q<350> q<351> q<352> q<353> q<354> 
+ q<355> q<356> q<357> q<358> q<359> q<360> q<361> q<362> q<363> q<364> q<365> 
+ q<366> q<367> q<368> q<369> q<370> q<371> q<372> q<373> q<374> q<375> q<376> 
+ q<377> q<378> q<379> q<380> q<381> q<382> q<383> q<384> q<385> q<386> q<387> 
+ q<388> q<389> q<390> q<391> q<392> q<393> q<394> q<395> q<396> q<397> q<398> 
+ q<399> q<400> q<401> q<402> q<403> q<404> q<405> q<406> q<407> q<408> q<409> 
+ q<410> q<411> q<412> q<413> q<414> q<415> q<416> q<417> q<418> q<419> q<420> 
+ q<421> q<422> q<423> q<424> q<425> q<426> q<427> q<428> q<429> q<430> q<431> 
+ q<432> q<433> q<434> q<435> q<436> q<437> q<438> q<439> q<440> q<441> q<442> 
+ q<443> q<444> q<445> q<446> q<447> q<448> q<449> q<450> q<451> q<452> q<453> 
+ q<454> q<455> q<456> q<457> q<458> q<459> q<460> q<461> q<462> q<463> q<464> 
+ q<465> q<466> q<467> q<468> q<469> q<470> q<471> q<472> q<473> q<474> q<475> 
+ q<476> q<477> q<478> q<479> q<480> q<481> q<482> q<483> q<484> q<485> q<486> 
+ q<487> q<488> q<489> q<490> q<491> q<492> q<493> q<494> q<495> q<496> q<497> 
+ q<498> q<499> q<500> q<501> q<502> q<503> q<504> q<505> q<506> q<507> q<508> 
+ q<509> q<510> q<511> time<0> time<1> time<2> time<3> vdd vss / 
+ Tgenerate_array_64
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    timegenerate
* View Name:    schematic
************************************************************************

.SUBCKT timegenerate entime in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> 
+ in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> 
+ in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> 
+ in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> 
+ in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> 
+ in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> 
+ in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> 
+ in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> 
+ in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> 
+ in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> 
+ in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> 
+ in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> 
+ in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> in1<113> 
+ in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> 
+ in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> in2<2> 
+ in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> 
+ in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> 
+ in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> 
+ in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> in2<39> 
+ in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> in2<48> 
+ in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> in2<57> 
+ in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> in2<66> 
+ in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> 
+ in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> in2<84> 
+ in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> 
+ in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> in2<102> 
+ in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> in2<110> 
+ in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> in2<118> 
+ in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> in2<126> 
+ in2<127> q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> 
+ q<13> q<14> q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> 
+ q<25> q<26> q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> 
+ q<37> q<38> q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> 
+ q<49> q<50> q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> 
+ q<61> q<62> q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> 
+ q<73> q<74> q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> 
+ q<85> q<86> q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> 
+ q<97> q<98> q<99> q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> 
+ q<108> q<109> q<110> q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> 
+ q<119> q<120> q<121> q<122> q<123> q<124> q<125> q<126> q<127> q<128> q<129> 
+ q<130> q<131> q<132> q<133> q<134> q<135> q<136> q<137> q<138> q<139> q<140> 
+ q<141> q<142> q<143> q<144> q<145> q<146> q<147> q<148> q<149> q<150> q<151> 
+ q<152> q<153> q<154> q<155> q<156> q<157> q<158> q<159> q<160> q<161> q<162> 
+ q<163> q<164> q<165> q<166> q<167> q<168> q<169> q<170> q<171> q<172> q<173> 
+ q<174> q<175> q<176> q<177> q<178> q<179> q<180> q<181> q<182> q<183> q<184> 
+ q<185> q<186> q<187> q<188> q<189> q<190> q<191> q<192> q<193> q<194> q<195> 
+ q<196> q<197> q<198> q<199> q<200> q<201> q<202> q<203> q<204> q<205> q<206> 
+ q<207> q<208> q<209> q<210> q<211> q<212> q<213> q<214> q<215> q<216> q<217> 
+ q<218> q<219> q<220> q<221> q<222> q<223> q<224> q<225> q<226> q<227> q<228> 
+ q<229> q<230> q<231> q<232> q<233> q<234> q<235> q<236> q<237> q<238> q<239> 
+ q<240> q<241> q<242> q<243> q<244> q<245> q<246> q<247> q<248> q<249> q<250> 
+ q<251> q<252> q<253> q<254> q<255> q<256> q<257> q<258> q<259> q<260> q<261> 
+ q<262> q<263> q<264> q<265> q<266> q<267> q<268> q<269> q<270> q<271> q<272> 
+ q<273> q<274> q<275> q<276> q<277> q<278> q<279> q<280> q<281> q<282> q<283> 
+ q<284> q<285> q<286> q<287> q<288> q<289> q<290> q<291> q<292> q<293> q<294> 
+ q<295> q<296> q<297> q<298> q<299> q<300> q<301> q<302> q<303> q<304> q<305> 
+ q<306> q<307> q<308> q<309> q<310> q<311> q<312> q<313> q<314> q<315> q<316> 
+ q<317> q<318> q<319> q<320> q<321> q<322> q<323> q<324> q<325> q<326> q<327> 
+ q<328> q<329> q<330> q<331> q<332> q<333> q<334> q<335> q<336> q<337> q<338> 
+ q<339> q<340> q<341> q<342> q<343> q<344> q<345> q<346> q<347> q<348> q<349> 
+ q<350> q<351> q<352> q<353> q<354> q<355> q<356> q<357> q<358> q<359> q<360> 
+ q<361> q<362> q<363> q<364> q<365> q<366> q<367> q<368> q<369> q<370> q<371> 
+ q<372> q<373> q<374> q<375> q<376> q<377> q<378> q<379> q<380> q<381> q<382> 
+ q<383> q<384> q<385> q<386> q<387> q<388> q<389> q<390> q<391> q<392> q<393> 
+ q<394> q<395> q<396> q<397> q<398> q<399> q<400> q<401> q<402> q<403> q<404> 
+ q<405> q<406> q<407> q<408> q<409> q<410> q<411> q<412> q<413> q<414> q<415> 
+ q<416> q<417> q<418> q<419> q<420> q<421> q<422> q<423> q<424> q<425> q<426> 
+ q<427> q<428> q<429> q<430> q<431> q<432> q<433> q<434> q<435> q<436> q<437> 
+ q<438> q<439> q<440> q<441> q<442> q<443> q<444> q<445> q<446> q<447> q<448> 
+ q<449> q<450> q<451> q<452> q<453> q<454> q<455> q<456> q<457> q<458> q<459> 
+ q<460> q<461> q<462> q<463> q<464> q<465> q<466> q<467> q<468> q<469> q<470> 
+ q<471> q<472> q<473> q<474> q<475> q<476> q<477> q<478> q<479> q<480> q<481> 
+ q<482> q<483> q<484> q<485> q<486> q<487> q<488> q<489> q<490> q<491> q<492> 
+ q<493> q<494> q<495> q<496> q<497> q<498> q<499> q<500> q<501> q<502> q<503> 
+ q<504> q<505> q<506> q<507> q<508> q<509> q<510> q<511> time<0> time<1> 
+ time<2> time<3> vdd vss
*.PININFO entime:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO q<16>:I q<17>:I q<18>:I q<19>:I q<20>:I q<21>:I q<22>:I q<23>:I 
*.PININFO q<24>:I q<25>:I q<26>:I q<27>:I q<28>:I q<29>:I q<30>:I q<31>:I 
*.PININFO q<32>:I q<33>:I q<34>:I q<35>:I q<36>:I q<37>:I q<38>:I q<39>:I 
*.PININFO q<40>:I q<41>:I q<42>:I q<43>:I q<44>:I q<45>:I q<46>:I q<47>:I 
*.PININFO q<48>:I q<49>:I q<50>:I q<51>:I q<52>:I q<53>:I q<54>:I q<55>:I 
*.PININFO q<56>:I q<57>:I q<58>:I q<59>:I q<60>:I q<61>:I q<62>:I q<63>:I 
*.PININFO q<64>:I q<65>:I q<66>:I q<67>:I q<68>:I q<69>:I q<70>:I q<71>:I 
*.PININFO q<72>:I q<73>:I q<74>:I q<75>:I q<76>:I q<77>:I q<78>:I q<79>:I 
*.PININFO q<80>:I q<81>:I q<82>:I q<83>:I q<84>:I q<85>:I q<86>:I q<87>:I 
*.PININFO q<88>:I q<89>:I q<90>:I q<91>:I q<92>:I q<93>:I q<94>:I q<95>:I 
*.PININFO q<96>:I q<97>:I q<98>:I q<99>:I q<100>:I q<101>:I q<102>:I q<103>:I 
*.PININFO q<104>:I q<105>:I q<106>:I q<107>:I q<108>:I q<109>:I q<110>:I 
*.PININFO q<111>:I q<112>:I q<113>:I q<114>:I q<115>:I q<116>:I q<117>:I 
*.PININFO q<118>:I q<119>:I q<120>:I q<121>:I q<122>:I q<123>:I q<124>:I 
*.PININFO q<125>:I q<126>:I q<127>:I q<128>:I q<129>:I q<130>:I q<131>:I 
*.PININFO q<132>:I q<133>:I q<134>:I q<135>:I q<136>:I q<137>:I q<138>:I 
*.PININFO q<139>:I q<140>:I q<141>:I q<142>:I q<143>:I q<144>:I q<145>:I 
*.PININFO q<146>:I q<147>:I q<148>:I q<149>:I q<150>:I q<151>:I q<152>:I 
*.PININFO q<153>:I q<154>:I q<155>:I q<156>:I q<157>:I q<158>:I q<159>:I 
*.PININFO q<160>:I q<161>:I q<162>:I q<163>:I q<164>:I q<165>:I q<166>:I 
*.PININFO q<167>:I q<168>:I q<169>:I q<170>:I q<171>:I q<172>:I q<173>:I 
*.PININFO q<174>:I q<175>:I q<176>:I q<177>:I q<178>:I q<179>:I q<180>:I 
*.PININFO q<181>:I q<182>:I q<183>:I q<184>:I q<185>:I q<186>:I q<187>:I 
*.PININFO q<188>:I q<189>:I q<190>:I q<191>:I q<192>:I q<193>:I q<194>:I 
*.PININFO q<195>:I q<196>:I q<197>:I q<198>:I q<199>:I q<200>:I q<201>:I 
*.PININFO q<202>:I q<203>:I q<204>:I q<205>:I q<206>:I q<207>:I q<208>:I 
*.PININFO q<209>:I q<210>:I q<211>:I q<212>:I q<213>:I q<214>:I q<215>:I 
*.PININFO q<216>:I q<217>:I q<218>:I q<219>:I q<220>:I q<221>:I q<222>:I 
*.PININFO q<223>:I q<224>:I q<225>:I q<226>:I q<227>:I q<228>:I q<229>:I 
*.PININFO q<230>:I q<231>:I q<232>:I q<233>:I q<234>:I q<235>:I q<236>:I 
*.PININFO q<237>:I q<238>:I q<239>:I q<240>:I q<241>:I q<242>:I q<243>:I 
*.PININFO q<244>:I q<245>:I q<246>:I q<247>:I q<248>:I q<249>:I q<250>:I 
*.PININFO q<251>:I q<252>:I q<253>:I q<254>:I q<255>:I q<256>:I q<257>:I 
*.PININFO q<258>:I q<259>:I q<260>:I q<261>:I q<262>:I q<263>:I q<264>:I 
*.PININFO q<265>:I q<266>:I q<267>:I q<268>:I q<269>:I q<270>:I q<271>:I 
*.PININFO q<272>:I q<273>:I q<274>:I q<275>:I q<276>:I q<277>:I q<278>:I 
*.PININFO q<279>:I q<280>:I q<281>:I q<282>:I q<283>:I q<284>:I q<285>:I 
*.PININFO q<286>:I q<287>:I q<288>:I q<289>:I q<290>:I q<291>:I q<292>:I 
*.PININFO q<293>:I q<294>:I q<295>:I q<296>:I q<297>:I q<298>:I q<299>:I 
*.PININFO q<300>:I q<301>:I q<302>:I q<303>:I q<304>:I q<305>:I q<306>:I 
*.PININFO q<307>:I q<308>:I q<309>:I q<310>:I q<311>:I q<312>:I q<313>:I 
*.PININFO q<314>:I q<315>:I q<316>:I q<317>:I q<318>:I q<319>:I q<320>:I 
*.PININFO q<321>:I q<322>:I q<323>:I q<324>:I q<325>:I q<326>:I q<327>:I 
*.PININFO q<328>:I q<329>:I q<330>:I q<331>:I q<332>:I q<333>:I q<334>:I 
*.PININFO q<335>:I q<336>:I q<337>:I q<338>:I q<339>:I q<340>:I q<341>:I 
*.PININFO q<342>:I q<343>:I q<344>:I q<345>:I q<346>:I q<347>:I q<348>:I 
*.PININFO q<349>:I q<350>:I q<351>:I q<352>:I q<353>:I q<354>:I q<355>:I 
*.PININFO q<356>:I q<357>:I q<358>:I q<359>:I q<360>:I q<361>:I q<362>:I 
*.PININFO q<363>:I q<364>:I q<365>:I q<366>:I q<367>:I q<368>:I q<369>:I 
*.PININFO q<370>:I q<371>:I q<372>:I q<373>:I q<374>:I q<375>:I q<376>:I 
*.PININFO q<377>:I q<378>:I q<379>:I q<380>:I q<381>:I q<382>:I q<383>:I 
*.PININFO q<384>:I q<385>:I q<386>:I q<387>:I q<388>:I q<389>:I q<390>:I 
*.PININFO q<391>:I q<392>:I q<393>:I q<394>:I q<395>:I q<396>:I q<397>:I 
*.PININFO q<398>:I q<399>:I q<400>:I q<401>:I q<402>:I q<403>:I q<404>:I 
*.PININFO q<405>:I q<406>:I q<407>:I q<408>:I q<409>:I q<410>:I q<411>:I 
*.PININFO q<412>:I q<413>:I q<414>:I q<415>:I q<416>:I q<417>:I q<418>:I 
*.PININFO q<419>:I q<420>:I q<421>:I q<422>:I q<423>:I q<424>:I q<425>:I 
*.PININFO q<426>:I q<427>:I q<428>:I q<429>:I q<430>:I q<431>:I q<432>:I 
*.PININFO q<433>:I q<434>:I q<435>:I q<436>:I q<437>:I q<438>:I q<439>:I 
*.PININFO q<440>:I q<441>:I q<442>:I q<443>:I q<444>:I q<445>:I q<446>:I 
*.PININFO q<447>:I q<448>:I q<449>:I q<450>:I q<451>:I q<452>:I q<453>:I 
*.PININFO q<454>:I q<455>:I q<456>:I q<457>:I q<458>:I q<459>:I q<460>:I 
*.PININFO q<461>:I q<462>:I q<463>:I q<464>:I q<465>:I q<466>:I q<467>:I 
*.PININFO q<468>:I q<469>:I q<470>:I q<471>:I q<472>:I q<473>:I q<474>:I 
*.PININFO q<475>:I q<476>:I q<477>:I q<478>:I q<479>:I q<480>:I q<481>:I 
*.PININFO q<482>:I q<483>:I q<484>:I q<485>:I q<486>:I q<487>:I q<488>:I 
*.PININFO q<489>:I q<490>:I q<491>:I q<492>:I q<493>:I q<494>:I q<495>:I 
*.PININFO q<496>:I q<497>:I q<498>:I q<499>:I q<500>:I q<501>:I q<502>:I 
*.PININFO q<503>:I q<504>:I q<505>:I q<506>:I q<507>:I q<508>:I q<509>:I 
*.PININFO q<510>:I q<511>:I time<0>:I time<1>:I time<2>:I time<3>:I in1<0>:O 
*.PININFO in1<1>:O in1<2>:O in1<3>:O in1<4>:O in1<5>:O in1<6>:O in1<7>:O 
*.PININFO in1<8>:O in1<9>:O in1<10>:O in1<11>:O in1<12>:O in1<13>:O in1<14>:O 
*.PININFO in1<15>:O in1<16>:O in1<17>:O in1<18>:O in1<19>:O in1<20>:O 
*.PININFO in1<21>:O in1<22>:O in1<23>:O in1<24>:O in1<25>:O in1<26>:O 
*.PININFO in1<27>:O in1<28>:O in1<29>:O in1<30>:O in1<31>:O in1<32>:O 
*.PININFO in1<33>:O in1<34>:O in1<35>:O in1<36>:O in1<37>:O in1<38>:O 
*.PININFO in1<39>:O in1<40>:O in1<41>:O in1<42>:O in1<43>:O in1<44>:O 
*.PININFO in1<45>:O in1<46>:O in1<47>:O in1<48>:O in1<49>:O in1<50>:O 
*.PININFO in1<51>:O in1<52>:O in1<53>:O in1<54>:O in1<55>:O in1<56>:O 
*.PININFO in1<57>:O in1<58>:O in1<59>:O in1<60>:O in1<61>:O in1<62>:O 
*.PININFO in1<63>:O in1<64>:O in1<65>:O in1<66>:O in1<67>:O in1<68>:O 
*.PININFO in1<69>:O in1<70>:O in1<71>:O in1<72>:O in1<73>:O in1<74>:O 
*.PININFO in1<75>:O in1<76>:O in1<77>:O in1<78>:O in1<79>:O in1<80>:O 
*.PININFO in1<81>:O in1<82>:O in1<83>:O in1<84>:O in1<85>:O in1<86>:O 
*.PININFO in1<87>:O in1<88>:O in1<89>:O in1<90>:O in1<91>:O in1<92>:O 
*.PININFO in1<93>:O in1<94>:O in1<95>:O in1<96>:O in1<97>:O in1<98>:O 
*.PININFO in1<99>:O in1<100>:O in1<101>:O in1<102>:O in1<103>:O in1<104>:O 
*.PININFO in1<105>:O in1<106>:O in1<107>:O in1<108>:O in1<109>:O in1<110>:O 
*.PININFO in1<111>:O in1<112>:O in1<113>:O in1<114>:O in1<115>:O in1<116>:O 
*.PININFO in1<117>:O in1<118>:O in1<119>:O in1<120>:O in1<121>:O in1<122>:O 
*.PININFO in1<123>:O in1<124>:O in1<125>:O in1<126>:O in1<127>:O in2<0>:O 
*.PININFO in2<1>:O in2<2>:O in2<3>:O in2<4>:O in2<5>:O in2<6>:O in2<7>:O 
*.PININFO in2<8>:O in2<9>:O in2<10>:O in2<11>:O in2<12>:O in2<13>:O in2<14>:O 
*.PININFO in2<15>:O in2<16>:O in2<17>:O in2<18>:O in2<19>:O in2<20>:O 
*.PININFO in2<21>:O in2<22>:O in2<23>:O in2<24>:O in2<25>:O in2<26>:O 
*.PININFO in2<27>:O in2<28>:O in2<29>:O in2<30>:O in2<31>:O in2<32>:O 
*.PININFO in2<33>:O in2<34>:O in2<35>:O in2<36>:O in2<37>:O in2<38>:O 
*.PININFO in2<39>:O in2<40>:O in2<41>:O in2<42>:O in2<43>:O in2<44>:O 
*.PININFO in2<45>:O in2<46>:O in2<47>:O in2<48>:O in2<49>:O in2<50>:O 
*.PININFO in2<51>:O in2<52>:O in2<53>:O in2<54>:O in2<55>:O in2<56>:O 
*.PININFO in2<57>:O in2<58>:O in2<59>:O in2<60>:O in2<61>:O in2<62>:O 
*.PININFO in2<63>:O in2<64>:O in2<65>:O in2<66>:O in2<67>:O in2<68>:O 
*.PININFO in2<69>:O in2<70>:O in2<71>:O in2<72>:O in2<73>:O in2<74>:O 
*.PININFO in2<75>:O in2<76>:O in2<77>:O in2<78>:O in2<79>:O in2<80>:O 
*.PININFO in2<81>:O in2<82>:O in2<83>:O in2<84>:O in2<85>:O in2<86>:O 
*.PININFO in2<87>:O in2<88>:O in2<89>:O in2<90>:O in2<91>:O in2<92>:O 
*.PININFO in2<93>:O in2<94>:O in2<95>:O in2<96>:O in2<97>:O in2<98>:O 
*.PININFO in2<99>:O in2<100>:O in2<101>:O in2<102>:O in2<103>:O in2<104>:O 
*.PININFO in2<105>:O in2<106>:O in2<107>:O in2<108>:O in2<109>:O in2<110>:O 
*.PININFO in2<111>:O in2<112>:O in2<113>:O in2<114>:O in2<115>:O in2<116>:O 
*.PININFO in2<117>:O in2<118>:O in2<119>:O in2<120>:O in2<121>:O in2<122>:O 
*.PININFO in2<123>:O in2<124>:O in2<125>:O in2<126>:O in2<127>:O vdd:B vss:B
XI10 entimeb in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> in1<8> 
+ in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> in1<17> 
+ in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> in1<26> 
+ in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> in1<35> 
+ in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> in1<44> 
+ in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> in1<53> 
+ in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> in1<62> 
+ in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> in1<71> 
+ in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> in1<80> 
+ in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> in1<89> 
+ in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> in1<98> 
+ in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> in1<106> 
+ in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> in1<113> in1<114> 
+ in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> in1<122> 
+ in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> in2<2> in2<3> 
+ in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> in2<13> 
+ in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> in2<22> 
+ in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> in2<31> 
+ in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> in2<39> in2<40> 
+ in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> in2<48> in2<49> 
+ in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> in2<57> in2<58> 
+ in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> in2<66> in2<67> 
+ in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> in2<76> 
+ in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> in2<84> in2<85> 
+ in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> in2<94> 
+ in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> in2<102> in2<103> 
+ in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> in2<110> in2<111> 
+ in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> in2<118> in2<119> 
+ in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> in2<126> in2<127> q<0> 
+ q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> 
+ q<15> q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> 
+ q<27> q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> q<37> q<38> 
+ q<39> q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> q<49> q<50> 
+ q<51> q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> q<61> q<62> 
+ q<63> q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> q<73> q<74> 
+ q<75> q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> q<85> q<86> 
+ q<87> q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> q<97> q<98> 
+ q<99> q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> q<108> q<109> 
+ q<110> q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> q<119> q<120> 
+ q<121> q<122> q<123> q<124> q<125> q<126> q<127> q<128> q<129> q<130> q<131> 
+ q<132> q<133> q<134> q<135> q<136> q<137> q<138> q<139> q<140> q<141> q<142> 
+ q<143> q<144> q<145> q<146> q<147> q<148> q<149> q<150> q<151> q<152> q<153> 
+ q<154> q<155> q<156> q<157> q<158> q<159> q<160> q<161> q<162> q<163> q<164> 
+ q<165> q<166> q<167> q<168> q<169> q<170> q<171> q<172> q<173> q<174> q<175> 
+ q<176> q<177> q<178> q<179> q<180> q<181> q<182> q<183> q<184> q<185> q<186> 
+ q<187> q<188> q<189> q<190> q<191> q<192> q<193> q<194> q<195> q<196> q<197> 
+ q<198> q<199> q<200> q<201> q<202> q<203> q<204> q<205> q<206> q<207> q<208> 
+ q<209> q<210> q<211> q<212> q<213> q<214> q<215> q<216> q<217> q<218> q<219> 
+ q<220> q<221> q<222> q<223> q<224> q<225> q<226> q<227> q<228> q<229> q<230> 
+ q<231> q<232> q<233> q<234> q<235> q<236> q<237> q<238> q<239> q<240> q<241> 
+ q<242> q<243> q<244> q<245> q<246> q<247> q<248> q<249> q<250> q<251> q<252> 
+ q<253> q<254> q<255> q<256> q<257> q<258> q<259> q<260> q<261> q<262> q<263> 
+ q<264> q<265> q<266> q<267> q<268> q<269> q<270> q<271> q<272> q<273> q<274> 
+ q<275> q<276> q<277> q<278> q<279> q<280> q<281> q<282> q<283> q<284> q<285> 
+ q<286> q<287> q<288> q<289> q<290> q<291> q<292> q<293> q<294> q<295> q<296> 
+ q<297> q<298> q<299> q<300> q<301> q<302> q<303> q<304> q<305> q<306> q<307> 
+ q<308> q<309> q<310> q<311> q<312> q<313> q<314> q<315> q<316> q<317> q<318> 
+ q<319> q<320> q<321> q<322> q<323> q<324> q<325> q<326> q<327> q<328> q<329> 
+ q<330> q<331> q<332> q<333> q<334> q<335> q<336> q<337> q<338> q<339> q<340> 
+ q<341> q<342> q<343> q<344> q<345> q<346> q<347> q<348> q<349> q<350> q<351> 
+ q<352> q<353> q<354> q<355> q<356> q<357> q<358> q<359> q<360> q<361> q<362> 
+ q<363> q<364> q<365> q<366> q<367> q<368> q<369> q<370> q<371> q<372> q<373> 
+ q<374> q<375> q<376> q<377> q<378> q<379> q<380> q<381> q<382> q<383> q<384> 
+ q<385> q<386> q<387> q<388> q<389> q<390> q<391> q<392> q<393> q<394> q<395> 
+ q<396> q<397> q<398> q<399> q<400> q<401> q<402> q<403> q<404> q<405> q<406> 
+ q<407> q<408> q<409> q<410> q<411> q<412> q<413> q<414> q<415> q<416> q<417> 
+ q<418> q<419> q<420> q<421> q<422> q<423> q<424> q<425> q<426> q<427> q<428> 
+ q<429> q<430> q<431> q<432> q<433> q<434> q<435> q<436> q<437> q<438> q<439> 
+ q<440> q<441> q<442> q<443> q<444> q<445> q<446> q<447> q<448> q<449> q<450> 
+ q<451> q<452> q<453> q<454> q<455> q<456> q<457> q<458> q<459> q<460> q<461> 
+ q<462> q<463> q<464> q<465> q<466> q<467> q<468> q<469> q<470> q<471> q<472> 
+ q<473> q<474> q<475> q<476> q<477> q<478> q<479> q<480> q<481> q<482> q<483> 
+ q<484> q<485> q<486> q<487> q<488> q<489> q<490> q<491> q<492> q<493> q<494> 
+ q<495> q<496> q<497> q<498> q<499> q<500> q<501> q<502> q<503> q<504> q<505> 
+ q<506> q<507> q<508> q<509> q<510> q<511> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate_array_128
XI2 net09 entimeb vdd vss / inv8
XI1<0> net019<0> timeb<0> vdd vss / inv8
XI1<1> net019<1> timeb<1> vdd vss / inv8
XI1<2> net019<2> timeb<2> vdd vss / inv8
XI1<3> net019<3> timeb<3> vdd vss / inv8
XI3 entime net09 vdd vss / inv4
XI25<0> time<0> net019<0> vdd vss / inv4
XI25<1> time<1> net019<1> vdd vss / inv4
XI25<2> time<2> net019<2> vdd vss / inv4
XI25<3> time<3> net019<3> vdd vss / inv4
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    mux8x1
* View Name:    schematic
************************************************************************

.SUBCKT mux8x1 group<0> group<1> group<2> group<3> group<4> group<5> group<6> 
+ group<7> in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> vdd vss
*.PININFO group<0>:I group<1>:I group<2>:I group<3>:I group<4>:I group<5>:I 
*.PININFO group<6>:I group<7>:I in:I out<0>:O out<1>:O out<2>:O out<3>:O 
*.PININFO out<4>:O out<5>:O out<6>:O out<7>:O vdd:B vss:B
XI19 net80 out<0> vdd vss / inv8
XI17 net81 out<1> vdd vss / inv8
XI6 net82 out<2> vdd vss / inv8
XI7 net83 out<3> vdd vss / inv8
XI9 net84 out<4> vdd vss / inv8
XI11 net85 out<5> vdd vss / inv8
XI13 net86 out<6> vdd vss / inv8
XI15 net87 out<7> vdd vss / inv8
XI23 in group<0> net80 vdd vss / nand
XI22 in group<1> net81 vdd vss / nand
XI21 in group<2> net82 vdd vss / nand
XI4 in group<7> net87 vdd vss / nand
XI0 in group<3> net83 vdd vss / nand
XI1 in group<4> net84 vdd vss / nand
XI2 in group<5> net85 vdd vss / nand
XI3 in group<6> net86 vdd vss / nand
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    WLdriver_editable
* View Name:    schematic
************************************************************************

.SUBCKT WLdriver_editable group<0> group<1> group<2> group<3> group<4> 
+ group<5> group<6> group<7> in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> 
+ in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> 
+ in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> 
+ in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> 
+ in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> 
+ in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> 
+ in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> 
+ in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> 
+ in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> 
+ in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> 
+ in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> 
+ in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> 
+ in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> in1<113> 
+ in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> 
+ in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> in2<2> 
+ in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> 
+ in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> 
+ in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> 
+ in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> in2<39> 
+ in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> in2<48> 
+ in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> in2<57> 
+ in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> in2<66> 
+ in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> 
+ in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> in2<84> 
+ in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> 
+ in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> in2<102> 
+ in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> in2<110> 
+ in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> in2<118> 
+ in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> in2<126> 
+ in2<127> row16<0> row16<1> row16<2> row16<3> row16<4> row16<5> row16<6> 
+ row16<7> row16<8> row16<9> row16<10> row16<11> row16<12> row16<13> row16<14> 
+ row16<15> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> 
+ wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> 
+ wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> 
+ wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> 
+ wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> 
+ wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> 
+ wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> 
+ wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> 
+ wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> 
+ wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127>
*.PININFO group<0>:I group<1>:I group<2>:I group<3>:I group<4>:I group<5>:I 
*.PININFO group<6>:I group<7>:I row16<0>:I row16<1>:I row16<2>:I row16<3>:I 
*.PININFO row16<4>:I row16<5>:I row16<6>:I row16<7>:I row16<8>:I row16<9>:I 
*.PININFO row16<10>:I row16<11>:I row16<12>:I row16<13>:I row16<14>:I 
*.PININFO row16<15>:I wl<0>:O wl<1>:O wl<2>:O wl<3>:O wl<4>:O wl<5>:O wl<6>:O 
*.PININFO wl<7>:O wl<8>:O wl<9>:O wl<10>:O wl<11>:O wl<12>:O wl<13>:O wl<14>:O 
*.PININFO wl<15>:O wl<16>:O wl<17>:O wl<18>:O wl<19>:O wl<20>:O wl<21>:O 
*.PININFO wl<22>:O wl<23>:O wl<24>:O wl<25>:O wl<26>:O wl<27>:O wl<28>:O 
*.PININFO wl<29>:O wl<30>:O wl<31>:O wl<32>:O wl<33>:O wl<34>:O wl<35>:O 
*.PININFO wl<36>:O wl<37>:O wl<38>:O wl<39>:O wl<40>:O wl<41>:O wl<42>:O 
*.PININFO wl<43>:O wl<44>:O wl<45>:O wl<46>:O wl<47>:O wl<48>:O wl<49>:O 
*.PININFO wl<50>:O wl<51>:O wl<52>:O wl<53>:O wl<54>:O wl<55>:O wl<56>:O 
*.PININFO wl<57>:O wl<58>:O wl<59>:O wl<60>:O wl<61>:O wl<62>:O wl<63>:O 
*.PININFO wl<64>:O wl<65>:O wl<66>:O wl<67>:O wl<68>:O wl<69>:O wl<70>:O 
*.PININFO wl<71>:O wl<72>:O wl<73>:O wl<74>:O wl<75>:O wl<76>:O wl<77>:O 
*.PININFO wl<78>:O wl<79>:O wl<80>:O wl<81>:O wl<82>:O wl<83>:O wl<84>:O 
*.PININFO wl<85>:O wl<86>:O wl<87>:O wl<88>:O wl<89>:O wl<90>:O wl<91>:O 
*.PININFO wl<92>:O wl<93>:O wl<94>:O wl<95>:O wl<96>:O wl<97>:O wl<98>:O 
*.PININFO wl<99>:O wl<100>:O wl<101>:O wl<102>:O wl<103>:O wl<104>:O wl<105>:O 
*.PININFO wl<106>:O wl<107>:O wl<108>:O wl<109>:O wl<110>:O wl<111>:O 
*.PININFO wl<112>:O wl<113>:O wl<114>:O wl<115>:O wl<116>:O wl<117>:O 
*.PININFO wl<118>:O wl<119>:O wl<120>:O wl<121>:O wl<122>:O wl<123>:O 
*.PININFO wl<124>:O wl<125>:O wl<126>:O wl<127>:O in1<0>:B in1<1>:B in1<2>:B 
*.PININFO in1<3>:B in1<4>:B in1<5>:B in1<6>:B in1<7>:B in1<8>:B in1<9>:B 
*.PININFO in1<10>:B in1<11>:B in1<12>:B in1<13>:B in1<14>:B in1<15>:B 
*.PININFO in1<16>:B in1<17>:B in1<18>:B in1<19>:B in1<20>:B in1<21>:B 
*.PININFO in1<22>:B in1<23>:B in1<24>:B in1<25>:B in1<26>:B in1<27>:B 
*.PININFO in1<28>:B in1<29>:B in1<30>:B in1<31>:B in1<32>:B in1<33>:B 
*.PININFO in1<34>:B in1<35>:B in1<36>:B in1<37>:B in1<38>:B in1<39>:B 
*.PININFO in1<40>:B in1<41>:B in1<42>:B in1<43>:B in1<44>:B in1<45>:B 
*.PININFO in1<46>:B in1<47>:B in1<48>:B in1<49>:B in1<50>:B in1<51>:B 
*.PININFO in1<52>:B in1<53>:B in1<54>:B in1<55>:B in1<56>:B in1<57>:B 
*.PININFO in1<58>:B in1<59>:B in1<60>:B in1<61>:B in1<62>:B in1<63>:B 
*.PININFO in1<64>:B in1<65>:B in1<66>:B in1<67>:B in1<68>:B in1<69>:B 
*.PININFO in1<70>:B in1<71>:B in1<72>:B in1<73>:B in1<74>:B in1<75>:B 
*.PININFO in1<76>:B in1<77>:B in1<78>:B in1<79>:B in1<80>:B in1<81>:B 
*.PININFO in1<82>:B in1<83>:B in1<84>:B in1<85>:B in1<86>:B in1<87>:B 
*.PININFO in1<88>:B in1<89>:B in1<90>:B in1<91>:B in1<92>:B in1<93>:B 
*.PININFO in1<94>:B in1<95>:B in1<96>:B in1<97>:B in1<98>:B in1<99>:B 
*.PININFO in1<100>:B in1<101>:B in1<102>:B in1<103>:B in1<104>:B in1<105>:B 
*.PININFO in1<106>:B in1<107>:B in1<108>:B in1<109>:B in1<110>:B in1<111>:B 
*.PININFO in1<112>:B in1<113>:B in1<114>:B in1<115>:B in1<116>:B in1<117>:B 
*.PININFO in1<118>:B in1<119>:B in1<120>:B in1<121>:B in1<122>:B in1<123>:B 
*.PININFO in1<124>:B in1<125>:B in1<126>:B in1<127>:B in2<0>:B in2<1>:B 
*.PININFO in2<2>:B in2<3>:B in2<4>:B in2<5>:B in2<6>:B in2<7>:B in2<8>:B 
*.PININFO in2<9>:B in2<10>:B in2<11>:B in2<12>:B in2<13>:B in2<14>:B in2<15>:B 
*.PININFO in2<16>:B in2<17>:B in2<18>:B in2<19>:B in2<20>:B in2<21>:B 
*.PININFO in2<22>:B in2<23>:B in2<24>:B in2<25>:B in2<26>:B in2<27>:B 
*.PININFO in2<28>:B in2<29>:B in2<30>:B in2<31>:B in2<32>:B in2<33>:B 
*.PININFO in2<34>:B in2<35>:B in2<36>:B in2<37>:B in2<38>:B in2<39>:B 
*.PININFO in2<40>:B in2<41>:B in2<42>:B in2<43>:B in2<44>:B in2<45>:B 
*.PININFO in2<46>:B in2<47>:B in2<48>:B in2<49>:B in2<50>:B in2<51>:B 
*.PININFO in2<52>:B in2<53>:B in2<54>:B in2<55>:B in2<56>:B in2<57>:B 
*.PININFO in2<58>:B in2<59>:B in2<60>:B in2<61>:B in2<62>:B in2<63>:B 
*.PININFO in2<64>:B in2<65>:B in2<66>:B in2<67>:B in2<68>:B in2<69>:B 
*.PININFO in2<70>:B in2<71>:B in2<72>:B in2<73>:B in2<74>:B in2<75>:B 
*.PININFO in2<76>:B in2<77>:B in2<78>:B in2<79>:B in2<80>:B in2<81>:B 
*.PININFO in2<82>:B in2<83>:B in2<84>:B in2<85>:B in2<86>:B in2<87>:B 
*.PININFO in2<88>:B in2<89>:B in2<90>:B in2<91>:B in2<92>:B in2<93>:B 
*.PININFO in2<94>:B in2<95>:B in2<96>:B in2<97>:B in2<98>:B in2<99>:B 
*.PININFO in2<100>:B in2<101>:B in2<102>:B in2<103>:B in2<104>:B in2<105>:B 
*.PININFO in2<106>:B in2<107>:B in2<108>:B in2<109>:B in2<110>:B in2<111>:B 
*.PININFO in2<112>:B in2<113>:B in2<114>:B in2<115>:B in2<116>:B in2<117>:B 
*.PININFO in2<118>:B in2<119>:B in2<120>:B in2<121>:B in2<122>:B in2<123>:B 
*.PININFO in2<124>:B in2<125>:B in2<126>:B in2<127>:B vdd:B vss:B
XI16 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<15> wl<120> wl<121> wl<122> wl<123> wl<124> wl<125> wl<126> wl<127> 
+ vdd vss / mux8x1
XI15 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<14> wl<112> wl<113> wl<114> wl<115> wl<116> wl<117> wl<118> wl<119> 
+ vdd vss / mux8x1
XI14 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<13> wl<104> wl<105> wl<106> wl<107> wl<108> wl<109> wl<110> wl<111> 
+ vdd vss / mux8x1
XI13 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<12> wl<96> wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> vdd 
+ vss / mux8x1
XI12 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<11> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> vdd vss / 
+ mux8x1
XI11 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<10> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> wl<86> wl<87> vdd vss / 
+ mux8x1
XI10 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<9> wl<72> wl<73> wl<74> wl<75> wl<76> wl<77> wl<78> wl<79> vdd vss / 
+ mux8x1
XI9 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<8> wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> vdd vss / 
+ mux8x1
XI8 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<7> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> vdd vss / 
+ mux8x1
XI7 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<6> wl<48> wl<49> wl<50> wl<51> wl<52> wl<53> wl<54> wl<55> vdd vss / 
+ mux8x1
XI6 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<5> wl<40> wl<41> wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> vdd vss / 
+ mux8x1
XI5 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<4> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> vdd vss / 
+ mux8x1
XI4 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<3> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> vdd vss / 
+ mux8x1
XI1 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<0> wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> vdd vss / mux8x1
XI2 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<1> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> vdd vss / 
+ mux8x1
XI3 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<2> wl<16> wl<17> wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> vdd vss / 
+ mux8x1
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    SRAMCIMfinal
* View Name:    schematic
************************************************************************

.SUBCKT SRAMCIMfinal a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> clk col_en comp 
+ d<31> d<30> d<29> d<28> d<27> d<26> d<25> d<24> d<23> d<22> d<21> d<20> 
+ d<19> d<18> d<17> d<16> d<15> d<14> d<13> d<12> d<11> d<10> d<9> d<8> d<7> 
+ d<6> d<5> d<4> d<3> d<2> d<1> d<0> data_in_cim<511> data_in_cim<510> 
+ data_in_cim<509> data_in_cim<508> data_in_cim<507> data_in_cim<506> 
+ data_in_cim<505> data_in_cim<504> data_in_cim<503> data_in_cim<502> 
+ data_in_cim<501> data_in_cim<500> data_in_cim<499> data_in_cim<498> 
+ data_in_cim<497> data_in_cim<496> data_in_cim<495> data_in_cim<494> 
+ data_in_cim<493> data_in_cim<492> data_in_cim<491> data_in_cim<490> 
+ data_in_cim<489> data_in_cim<488> data_in_cim<487> data_in_cim<486> 
+ data_in_cim<485> data_in_cim<484> data_in_cim<483> data_in_cim<482> 
+ data_in_cim<481> data_in_cim<480> data_in_cim<479> data_in_cim<478> 
+ data_in_cim<477> data_in_cim<476> data_in_cim<475> data_in_cim<474> 
+ data_in_cim<473> data_in_cim<472> data_in_cim<471> data_in_cim<470> 
+ data_in_cim<469> data_in_cim<468> data_in_cim<467> data_in_cim<466> 
+ data_in_cim<465> data_in_cim<464> data_in_cim<463> data_in_cim<462> 
+ data_in_cim<461> data_in_cim<460> data_in_cim<459> data_in_cim<458> 
+ data_in_cim<457> data_in_cim<456> data_in_cim<455> data_in_cim<454> 
+ data_in_cim<453> data_in_cim<452> data_in_cim<451> data_in_cim<450> 
+ data_in_cim<449> data_in_cim<448> data_in_cim<447> data_in_cim<446> 
+ data_in_cim<445> data_in_cim<444> data_in_cim<443> data_in_cim<442> 
+ data_in_cim<441> data_in_cim<440> data_in_cim<439> data_in_cim<438> 
+ data_in_cim<437> data_in_cim<436> data_in_cim<435> data_in_cim<434> 
+ data_in_cim<433> data_in_cim<432> data_in_cim<431> data_in_cim<430> 
+ data_in_cim<429> data_in_cim<428> data_in_cim<427> data_in_cim<426> 
+ data_in_cim<425> data_in_cim<424> data_in_cim<423> data_in_cim<422> 
+ data_in_cim<421> data_in_cim<420> data_in_cim<419> data_in_cim<418> 
+ data_in_cim<417> data_in_cim<416> data_in_cim<415> data_in_cim<414> 
+ data_in_cim<413> data_in_cim<412> data_in_cim<411> data_in_cim<410> 
+ data_in_cim<409> data_in_cim<408> data_in_cim<407> data_in_cim<406> 
+ data_in_cim<405> data_in_cim<404> data_in_cim<403> data_in_cim<402> 
+ data_in_cim<401> data_in_cim<400> data_in_cim<399> data_in_cim<398> 
+ data_in_cim<397> data_in_cim<396> data_in_cim<395> data_in_cim<394> 
+ data_in_cim<393> data_in_cim<392> data_in_cim<391> data_in_cim<390> 
+ data_in_cim<389> data_in_cim<388> data_in_cim<387> data_in_cim<386> 
+ data_in_cim<385> data_in_cim<384> data_in_cim<383> data_in_cim<382> 
+ data_in_cim<381> data_in_cim<380> data_in_cim<379> data_in_cim<378> 
+ data_in_cim<377> data_in_cim<376> data_in_cim<375> data_in_cim<374> 
+ data_in_cim<373> data_in_cim<372> data_in_cim<371> data_in_cim<370> 
+ data_in_cim<369> data_in_cim<368> data_in_cim<367> data_in_cim<366> 
+ data_in_cim<365> data_in_cim<364> data_in_cim<363> data_in_cim<362> 
+ data_in_cim<361> data_in_cim<360> data_in_cim<359> data_in_cim<358> 
+ data_in_cim<357> data_in_cim<356> data_in_cim<355> data_in_cim<354> 
+ data_in_cim<353> data_in_cim<352> data_in_cim<351> data_in_cim<350> 
+ data_in_cim<349> data_in_cim<348> data_in_cim<347> data_in_cim<346> 
+ data_in_cim<345> data_in_cim<344> data_in_cim<343> data_in_cim<342> 
+ data_in_cim<341> data_in_cim<340> data_in_cim<339> data_in_cim<338> 
+ data_in_cim<337> data_in_cim<336> data_in_cim<335> data_in_cim<334> 
+ data_in_cim<333> data_in_cim<332> data_in_cim<331> data_in_cim<330> 
+ data_in_cim<329> data_in_cim<328> data_in_cim<327> data_in_cim<326> 
+ data_in_cim<325> data_in_cim<324> data_in_cim<323> data_in_cim<322> 
+ data_in_cim<321> data_in_cim<320> data_in_cim<319> data_in_cim<318> 
+ data_in_cim<317> data_in_cim<316> data_in_cim<315> data_in_cim<314> 
+ data_in_cim<313> data_in_cim<312> data_in_cim<311> data_in_cim<310> 
+ data_in_cim<309> data_in_cim<308> data_in_cim<307> data_in_cim<306> 
+ data_in_cim<305> data_in_cim<304> data_in_cim<303> data_in_cim<302> 
+ data_in_cim<301> data_in_cim<300> data_in_cim<299> data_in_cim<298> 
+ data_in_cim<297> data_in_cim<296> data_in_cim<295> data_in_cim<294> 
+ data_in_cim<293> data_in_cim<292> data_in_cim<291> data_in_cim<290> 
+ data_in_cim<289> data_in_cim<288> data_in_cim<287> data_in_cim<286> 
+ data_in_cim<285> data_in_cim<284> data_in_cim<283> data_in_cim<282> 
+ data_in_cim<281> data_in_cim<280> data_in_cim<279> data_in_cim<278> 
+ data_in_cim<277> data_in_cim<276> data_in_cim<275> data_in_cim<274> 
+ data_in_cim<273> data_in_cim<272> data_in_cim<271> data_in_cim<270> 
+ data_in_cim<269> data_in_cim<268> data_in_cim<267> data_in_cim<266> 
+ data_in_cim<265> data_in_cim<264> data_in_cim<263> data_in_cim<262> 
+ data_in_cim<261> data_in_cim<260> data_in_cim<259> data_in_cim<258> 
+ data_in_cim<257> data_in_cim<256> data_in_cim<255> data_in_cim<254> 
+ data_in_cim<253> data_in_cim<252> data_in_cim<251> data_in_cim<250> 
+ data_in_cim<249> data_in_cim<248> data_in_cim<247> data_in_cim<246> 
+ data_in_cim<245> data_in_cim<244> data_in_cim<243> data_in_cim<242> 
+ data_in_cim<241> data_in_cim<240> data_in_cim<239> data_in_cim<238> 
+ data_in_cim<237> data_in_cim<236> data_in_cim<235> data_in_cim<234> 
+ data_in_cim<233> data_in_cim<232> data_in_cim<231> data_in_cim<230> 
+ data_in_cim<229> data_in_cim<228> data_in_cim<227> data_in_cim<226> 
+ data_in_cim<225> data_in_cim<224> data_in_cim<223> data_in_cim<222> 
+ data_in_cim<221> data_in_cim<220> data_in_cim<219> data_in_cim<218> 
+ data_in_cim<217> data_in_cim<216> data_in_cim<215> data_in_cim<214> 
+ data_in_cim<213> data_in_cim<212> data_in_cim<211> data_in_cim<210> 
+ data_in_cim<209> data_in_cim<208> data_in_cim<207> data_in_cim<206> 
+ data_in_cim<205> data_in_cim<204> data_in_cim<203> data_in_cim<202> 
+ data_in_cim<201> data_in_cim<200> data_in_cim<199> data_in_cim<198> 
+ data_in_cim<197> data_in_cim<196> data_in_cim<195> data_in_cim<194> 
+ data_in_cim<193> data_in_cim<192> data_in_cim<191> data_in_cim<190> 
+ data_in_cim<189> data_in_cim<188> data_in_cim<187> data_in_cim<186> 
+ data_in_cim<185> data_in_cim<184> data_in_cim<183> data_in_cim<182> 
+ data_in_cim<181> data_in_cim<180> data_in_cim<179> data_in_cim<178> 
+ data_in_cim<177> data_in_cim<176> data_in_cim<175> data_in_cim<174> 
+ data_in_cim<173> data_in_cim<172> data_in_cim<171> data_in_cim<170> 
+ data_in_cim<169> data_in_cim<168> data_in_cim<167> data_in_cim<166> 
+ data_in_cim<165> data_in_cim<164> data_in_cim<163> data_in_cim<162> 
+ data_in_cim<161> data_in_cim<160> data_in_cim<159> data_in_cim<158> 
+ data_in_cim<157> data_in_cim<156> data_in_cim<155> data_in_cim<154> 
+ data_in_cim<153> data_in_cim<152> data_in_cim<151> data_in_cim<150> 
+ data_in_cim<149> data_in_cim<148> data_in_cim<147> data_in_cim<146> 
+ data_in_cim<145> data_in_cim<144> data_in_cim<143> data_in_cim<142> 
+ data_in_cim<141> data_in_cim<140> data_in_cim<139> data_in_cim<138> 
+ data_in_cim<137> data_in_cim<136> data_in_cim<135> data_in_cim<134> 
+ data_in_cim<133> data_in_cim<132> data_in_cim<131> data_in_cim<130> 
+ data_in_cim<129> data_in_cim<128> data_in_cim<127> data_in_cim<126> 
+ data_in_cim<125> data_in_cim<124> data_in_cim<123> data_in_cim<122> 
+ data_in_cim<121> data_in_cim<120> data_in_cim<119> data_in_cim<118> 
+ data_in_cim<117> data_in_cim<116> data_in_cim<115> data_in_cim<114> 
+ data_in_cim<113> data_in_cim<112> data_in_cim<111> data_in_cim<110> 
+ data_in_cim<109> data_in_cim<108> data_in_cim<107> data_in_cim<106> 
+ data_in_cim<105> data_in_cim<104> data_in_cim<103> data_in_cim<102> 
+ data_in_cim<101> data_in_cim<100> data_in_cim<99> data_in_cim<98> 
+ data_in_cim<97> data_in_cim<96> data_in_cim<95> data_in_cim<94> 
+ data_in_cim<93> data_in_cim<92> data_in_cim<91> data_in_cim<90> 
+ data_in_cim<89> data_in_cim<88> data_in_cim<87> data_in_cim<86> 
+ data_in_cim<85> data_in_cim<84> data_in_cim<83> data_in_cim<82> 
+ data_in_cim<81> data_in_cim<80> data_in_cim<79> data_in_cim<78> 
+ data_in_cim<77> data_in_cim<76> data_in_cim<75> data_in_cim<74> 
+ data_in_cim<73> data_in_cim<72> data_in_cim<71> data_in_cim<70> 
+ data_in_cim<69> data_in_cim<68> data_in_cim<67> data_in_cim<66> 
+ data_in_cim<65> data_in_cim<64> data_in_cim<63> data_in_cim<62> 
+ data_in_cim<61> data_in_cim<60> data_in_cim<59> data_in_cim<58> 
+ data_in_cim<57> data_in_cim<56> data_in_cim<55> data_in_cim<54> 
+ data_in_cim<53> data_in_cim<52> data_in_cim<51> data_in_cim<50> 
+ data_in_cim<49> data_in_cim<48> data_in_cim<47> data_in_cim<46> 
+ data_in_cim<45> data_in_cim<44> data_in_cim<43> data_in_cim<42> 
+ data_in_cim<41> data_in_cim<40> data_in_cim<39> data_in_cim<38> 
+ data_in_cim<37> data_in_cim<36> data_in_cim<35> data_in_cim<34> 
+ data_in_cim<33> data_in_cim<32> data_in_cim<31> data_in_cim<30> 
+ data_in_cim<29> data_in_cim<28> data_in_cim<27> data_in_cim<26> 
+ data_in_cim<25> data_in_cim<24> data_in_cim<23> data_in_cim<22> 
+ data_in_cim<21> data_in_cim<20> data_in_cim<19> data_in_cim<18> 
+ data_in_cim<17> data_in_cim<16> data_in_cim<15> data_in_cim<14> 
+ data_in_cim<13> data_in_cim<12> data_in_cim<11> data_in_cim<10> 
+ data_in_cim<9> data_in_cim<8> data_in_cim<7> data_in_cim<6> data_in_cim<5> 
+ data_in_cim<4> data_in_cim<3> data_in_cim<2> data_in_cim<1> data_in_cim<0> 
+ inbit model q<191> q<190> q<189> q<188> q<187> q<186> q<185> q<184> q<183> 
+ q<182> q<181> q<180> q<179> q<178> q<177> q<176> q<175> q<174> q<173> q<172> 
+ q<171> q<170> q<169> q<168> q<167> q<166> q<165> q<164> q<163> q<162> q<161> 
+ q<160> q<159> q<158> q<157> q<156> q<155> q<154> q<153> q<152> q<151> q<150> 
+ q<149> q<148> q<147> q<146> q<145> q<144> q<143> q<142> q<141> q<140> q<139> 
+ q<138> q<137> q<136> q<135> q<134> q<133> q<132> q<131> q<130> q<129> q<128> 
+ q<127> q<126> q<125> q<124> q<123> q<122> q<121> q<120> q<119> q<118> q<117> 
+ q<116> q<115> q<114> q<113> q<112> q<111> q<110> q<109> q<108> q<107> q<106> 
+ q<105> q<104> q<103> q<102> q<101> q<100> q<99> q<98> q<97> q<96> q<95> 
+ q<94> q<93> q<92> q<91> q<90> q<89> q<88> q<87> q<86> q<85> q<84> q<83> 
+ q<82> q<81> q<80> q<79> q<78> q<77> q<76> q<75> q<74> q<73> q<72> q<71> 
+ q<70> q<69> q<68> q<67> q<66> q<65> q<64> q<63> q<62> q<61> q<60> q<59> 
+ q<58> q<57> q<56> q<55> q<54> q<53> q<52> q<51> q<50> q<49> q<48> q<47> 
+ q<46> q<45> q<44> q<43> q<42> q<41> q<40> q<39> q<38> q<37> q<36> q<35> 
+ q<34> q<33> q<32> q<31> q<30> q<29> q<28> q<27> q<26> q<25> q<24> q<23> 
+ q<22> q<21> q<20> q<19> q<18> q<17> q<16> q<15> q<14> q<13> q<12> q<11> 
+ q<10> q<9> q<8> q<7> q<6> q<5> q<4> q<3> q<2> q<1> q<0> reg_en sel_array<15> 
+ sel_array<14> sel_array<13> sel_array<12> sel_array<11> sel_array<10> 
+ sel_array<9> sel_array<8> sel_array<7> sel_array<6> sel_array<5> 
+ sel_array<4> sel_array<3> sel_array<2> sel_array<1> sel_array<0> set vdd vss 
+ wait_ wrt
*.PININFO a<7>:I a<6>:I a<5>:I a<4>:I a<3>:I a<2>:I a<1>:I a<0>:I clk:I 
*.PININFO col_en:I comp:I d<31>:I d<30>:I d<29>:I d<28>:I d<27>:I d<26>:I 
*.PININFO d<25>:I d<24>:I d<23>:I d<22>:I d<21>:I d<20>:I d<19>:I d<18>:I 
*.PININFO d<17>:I d<16>:I d<15>:I d<14>:I d<13>:I d<12>:I d<11>:I d<10>:I 
*.PININFO d<9>:I d<8>:I d<7>:I d<6>:I d<5>:I d<4>:I d<3>:I d<2>:I d<1>:I 
*.PININFO d<0>:I data_in_cim<511>:I data_in_cim<510>:I data_in_cim<509>:I 
*.PININFO data_in_cim<508>:I data_in_cim<507>:I data_in_cim<506>:I 
*.PININFO data_in_cim<505>:I data_in_cim<504>:I data_in_cim<503>:I 
*.PININFO data_in_cim<502>:I data_in_cim<501>:I data_in_cim<500>:I 
*.PININFO data_in_cim<499>:I data_in_cim<498>:I data_in_cim<497>:I 
*.PININFO data_in_cim<496>:I data_in_cim<495>:I data_in_cim<494>:I 
*.PININFO data_in_cim<493>:I data_in_cim<492>:I data_in_cim<491>:I 
*.PININFO data_in_cim<490>:I data_in_cim<489>:I data_in_cim<488>:I 
*.PININFO data_in_cim<487>:I data_in_cim<486>:I data_in_cim<485>:I 
*.PININFO data_in_cim<484>:I data_in_cim<483>:I data_in_cim<482>:I 
*.PININFO data_in_cim<481>:I data_in_cim<480>:I data_in_cim<479>:I 
*.PININFO data_in_cim<478>:I data_in_cim<477>:I data_in_cim<476>:I 
*.PININFO data_in_cim<475>:I data_in_cim<474>:I data_in_cim<473>:I 
*.PININFO data_in_cim<472>:I data_in_cim<471>:I data_in_cim<470>:I 
*.PININFO data_in_cim<469>:I data_in_cim<468>:I data_in_cim<467>:I 
*.PININFO data_in_cim<466>:I data_in_cim<465>:I data_in_cim<464>:I 
*.PININFO data_in_cim<463>:I data_in_cim<462>:I data_in_cim<461>:I 
*.PININFO data_in_cim<460>:I data_in_cim<459>:I data_in_cim<458>:I 
*.PININFO data_in_cim<457>:I data_in_cim<456>:I data_in_cim<455>:I 
*.PININFO data_in_cim<454>:I data_in_cim<453>:I data_in_cim<452>:I 
*.PININFO data_in_cim<451>:I data_in_cim<450>:I data_in_cim<449>:I 
*.PININFO data_in_cim<448>:I data_in_cim<447>:I data_in_cim<446>:I 
*.PININFO data_in_cim<445>:I data_in_cim<444>:I data_in_cim<443>:I 
*.PININFO data_in_cim<442>:I data_in_cim<441>:I data_in_cim<440>:I 
*.PININFO data_in_cim<439>:I data_in_cim<438>:I data_in_cim<437>:I 
*.PININFO data_in_cim<436>:I data_in_cim<435>:I data_in_cim<434>:I 
*.PININFO data_in_cim<433>:I data_in_cim<432>:I data_in_cim<431>:I 
*.PININFO data_in_cim<430>:I data_in_cim<429>:I data_in_cim<428>:I 
*.PININFO data_in_cim<427>:I data_in_cim<426>:I data_in_cim<425>:I 
*.PININFO data_in_cim<424>:I data_in_cim<423>:I data_in_cim<422>:I 
*.PININFO data_in_cim<421>:I data_in_cim<420>:I data_in_cim<419>:I 
*.PININFO data_in_cim<418>:I data_in_cim<417>:I data_in_cim<416>:I 
*.PININFO data_in_cim<415>:I data_in_cim<414>:I data_in_cim<413>:I 
*.PININFO data_in_cim<412>:I data_in_cim<411>:I data_in_cim<410>:I 
*.PININFO data_in_cim<409>:I data_in_cim<408>:I data_in_cim<407>:I 
*.PININFO data_in_cim<406>:I data_in_cim<405>:I data_in_cim<404>:I 
*.PININFO data_in_cim<403>:I data_in_cim<402>:I data_in_cim<401>:I 
*.PININFO data_in_cim<400>:I data_in_cim<399>:I data_in_cim<398>:I 
*.PININFO data_in_cim<397>:I data_in_cim<396>:I data_in_cim<395>:I 
*.PININFO data_in_cim<394>:I data_in_cim<393>:I data_in_cim<392>:I 
*.PININFO data_in_cim<391>:I data_in_cim<390>:I data_in_cim<389>:I 
*.PININFO data_in_cim<388>:I data_in_cim<387>:I data_in_cim<386>:I 
*.PININFO data_in_cim<385>:I data_in_cim<384>:I data_in_cim<383>:I 
*.PININFO data_in_cim<382>:I data_in_cim<381>:I data_in_cim<380>:I 
*.PININFO data_in_cim<379>:I data_in_cim<378>:I data_in_cim<377>:I 
*.PININFO data_in_cim<376>:I data_in_cim<375>:I data_in_cim<374>:I 
*.PININFO data_in_cim<373>:I data_in_cim<372>:I data_in_cim<371>:I 
*.PININFO data_in_cim<370>:I data_in_cim<369>:I data_in_cim<368>:I 
*.PININFO data_in_cim<367>:I data_in_cim<366>:I data_in_cim<365>:I 
*.PININFO data_in_cim<364>:I data_in_cim<363>:I data_in_cim<362>:I 
*.PININFO data_in_cim<361>:I data_in_cim<360>:I data_in_cim<359>:I 
*.PININFO data_in_cim<358>:I data_in_cim<357>:I data_in_cim<356>:I 
*.PININFO data_in_cim<355>:I data_in_cim<354>:I data_in_cim<353>:I 
*.PININFO data_in_cim<352>:I data_in_cim<351>:I data_in_cim<350>:I 
*.PININFO data_in_cim<349>:I data_in_cim<348>:I data_in_cim<347>:I 
*.PININFO data_in_cim<346>:I data_in_cim<345>:I data_in_cim<344>:I 
*.PININFO data_in_cim<343>:I data_in_cim<342>:I data_in_cim<341>:I 
*.PININFO data_in_cim<340>:I data_in_cim<339>:I data_in_cim<338>:I 
*.PININFO data_in_cim<337>:I data_in_cim<336>:I data_in_cim<335>:I 
*.PININFO data_in_cim<334>:I data_in_cim<333>:I data_in_cim<332>:I 
*.PININFO data_in_cim<331>:I data_in_cim<330>:I data_in_cim<329>:I 
*.PININFO data_in_cim<328>:I data_in_cim<327>:I data_in_cim<326>:I 
*.PININFO data_in_cim<325>:I data_in_cim<324>:I data_in_cim<323>:I 
*.PININFO data_in_cim<322>:I data_in_cim<321>:I data_in_cim<320>:I 
*.PININFO data_in_cim<319>:I data_in_cim<318>:I data_in_cim<317>:I 
*.PININFO data_in_cim<316>:I data_in_cim<315>:I data_in_cim<314>:I 
*.PININFO data_in_cim<313>:I data_in_cim<312>:I data_in_cim<311>:I 
*.PININFO data_in_cim<310>:I data_in_cim<309>:I data_in_cim<308>:I 
*.PININFO data_in_cim<307>:I data_in_cim<306>:I data_in_cim<305>:I 
*.PININFO data_in_cim<304>:I data_in_cim<303>:I data_in_cim<302>:I 
*.PININFO data_in_cim<301>:I data_in_cim<300>:I data_in_cim<299>:I 
*.PININFO data_in_cim<298>:I data_in_cim<297>:I data_in_cim<296>:I 
*.PININFO data_in_cim<295>:I data_in_cim<294>:I data_in_cim<293>:I 
*.PININFO data_in_cim<292>:I data_in_cim<291>:I data_in_cim<290>:I 
*.PININFO data_in_cim<289>:I data_in_cim<288>:I data_in_cim<287>:I 
*.PININFO data_in_cim<286>:I data_in_cim<285>:I data_in_cim<284>:I 
*.PININFO data_in_cim<283>:I data_in_cim<282>:I data_in_cim<281>:I 
*.PININFO data_in_cim<280>:I data_in_cim<279>:I data_in_cim<278>:I 
*.PININFO data_in_cim<277>:I data_in_cim<276>:I data_in_cim<275>:I 
*.PININFO data_in_cim<274>:I data_in_cim<273>:I data_in_cim<272>:I 
*.PININFO data_in_cim<271>:I data_in_cim<270>:I data_in_cim<269>:I 
*.PININFO data_in_cim<268>:I data_in_cim<267>:I data_in_cim<266>:I 
*.PININFO data_in_cim<265>:I data_in_cim<264>:I data_in_cim<263>:I 
*.PININFO data_in_cim<262>:I data_in_cim<261>:I data_in_cim<260>:I 
*.PININFO data_in_cim<259>:I data_in_cim<258>:I data_in_cim<257>:I 
*.PININFO data_in_cim<256>:I data_in_cim<255>:I data_in_cim<254>:I 
*.PININFO data_in_cim<253>:I data_in_cim<252>:I data_in_cim<251>:I 
*.PININFO data_in_cim<250>:I data_in_cim<249>:I data_in_cim<248>:I 
*.PININFO data_in_cim<247>:I data_in_cim<246>:I data_in_cim<245>:I 
*.PININFO data_in_cim<244>:I data_in_cim<243>:I data_in_cim<242>:I 
*.PININFO data_in_cim<241>:I data_in_cim<240>:I data_in_cim<239>:I 
*.PININFO data_in_cim<238>:I data_in_cim<237>:I data_in_cim<236>:I 
*.PININFO data_in_cim<235>:I data_in_cim<234>:I data_in_cim<233>:I 
*.PININFO data_in_cim<232>:I data_in_cim<231>:I data_in_cim<230>:I 
*.PININFO data_in_cim<229>:I data_in_cim<228>:I data_in_cim<227>:I 
*.PININFO data_in_cim<226>:I data_in_cim<225>:I data_in_cim<224>:I 
*.PININFO data_in_cim<223>:I data_in_cim<222>:I data_in_cim<221>:I 
*.PININFO data_in_cim<220>:I data_in_cim<219>:I data_in_cim<218>:I 
*.PININFO data_in_cim<217>:I data_in_cim<216>:I data_in_cim<215>:I 
*.PININFO data_in_cim<214>:I data_in_cim<213>:I data_in_cim<212>:I 
*.PININFO data_in_cim<211>:I data_in_cim<210>:I data_in_cim<209>:I 
*.PININFO data_in_cim<208>:I data_in_cim<207>:I data_in_cim<206>:I 
*.PININFO data_in_cim<205>:I data_in_cim<204>:I data_in_cim<203>:I 
*.PININFO data_in_cim<202>:I data_in_cim<201>:I data_in_cim<200>:I 
*.PININFO data_in_cim<199>:I data_in_cim<198>:I data_in_cim<197>:I 
*.PININFO data_in_cim<196>:I data_in_cim<195>:I data_in_cim<194>:I 
*.PININFO data_in_cim<193>:I data_in_cim<192>:I data_in_cim<191>:I 
*.PININFO data_in_cim<190>:I data_in_cim<189>:I data_in_cim<188>:I 
*.PININFO data_in_cim<187>:I data_in_cim<186>:I data_in_cim<185>:I 
*.PININFO data_in_cim<184>:I data_in_cim<183>:I data_in_cim<182>:I 
*.PININFO data_in_cim<181>:I data_in_cim<180>:I data_in_cim<179>:I 
*.PININFO data_in_cim<178>:I data_in_cim<177>:I data_in_cim<176>:I 
*.PININFO data_in_cim<175>:I data_in_cim<174>:I data_in_cim<173>:I 
*.PININFO data_in_cim<172>:I data_in_cim<171>:I data_in_cim<170>:I 
*.PININFO data_in_cim<169>:I data_in_cim<168>:I data_in_cim<167>:I 
*.PININFO data_in_cim<166>:I data_in_cim<165>:I data_in_cim<164>:I 
*.PININFO data_in_cim<163>:I data_in_cim<162>:I data_in_cim<161>:I 
*.PININFO data_in_cim<160>:I data_in_cim<159>:I data_in_cim<158>:I 
*.PININFO data_in_cim<157>:I data_in_cim<156>:I data_in_cim<155>:I 
*.PININFO data_in_cim<154>:I data_in_cim<153>:I data_in_cim<152>:I 
*.PININFO data_in_cim<151>:I data_in_cim<150>:I data_in_cim<149>:I 
*.PININFO data_in_cim<148>:I data_in_cim<147>:I data_in_cim<146>:I 
*.PININFO data_in_cim<145>:I data_in_cim<144>:I data_in_cim<143>:I 
*.PININFO data_in_cim<142>:I data_in_cim<141>:I data_in_cim<140>:I 
*.PININFO data_in_cim<139>:I data_in_cim<138>:I data_in_cim<137>:I 
*.PININFO data_in_cim<136>:I data_in_cim<135>:I data_in_cim<134>:I 
*.PININFO data_in_cim<133>:I data_in_cim<132>:I data_in_cim<131>:I 
*.PININFO data_in_cim<130>:I data_in_cim<129>:I data_in_cim<128>:I 
*.PININFO data_in_cim<127>:I data_in_cim<126>:I data_in_cim<125>:I 
*.PININFO data_in_cim<124>:I data_in_cim<123>:I data_in_cim<122>:I 
*.PININFO data_in_cim<121>:I data_in_cim<120>:I data_in_cim<119>:I 
*.PININFO data_in_cim<118>:I data_in_cim<117>:I data_in_cim<116>:I 
*.PININFO data_in_cim<115>:I data_in_cim<114>:I data_in_cim<113>:I 
*.PININFO data_in_cim<112>:I data_in_cim<111>:I data_in_cim<110>:I 
*.PININFO data_in_cim<109>:I data_in_cim<108>:I data_in_cim<107>:I 
*.PININFO data_in_cim<106>:I data_in_cim<105>:I data_in_cim<104>:I 
*.PININFO data_in_cim<103>:I data_in_cim<102>:I data_in_cim<101>:I 
*.PININFO data_in_cim<100>:I data_in_cim<99>:I data_in_cim<98>:I 
*.PININFO data_in_cim<97>:I data_in_cim<96>:I data_in_cim<95>:I 
*.PININFO data_in_cim<94>:I data_in_cim<93>:I data_in_cim<92>:I 
*.PININFO data_in_cim<91>:I data_in_cim<90>:I data_in_cim<89>:I 
*.PININFO data_in_cim<88>:I data_in_cim<87>:I data_in_cim<86>:I 
*.PININFO data_in_cim<85>:I data_in_cim<84>:I data_in_cim<83>:I 
*.PININFO data_in_cim<82>:I data_in_cim<81>:I data_in_cim<80>:I 
*.PININFO data_in_cim<79>:I data_in_cim<78>:I data_in_cim<77>:I 
*.PININFO data_in_cim<76>:I data_in_cim<75>:I data_in_cim<74>:I 
*.PININFO data_in_cim<73>:I data_in_cim<72>:I data_in_cim<71>:I 
*.PININFO data_in_cim<70>:I data_in_cim<69>:I data_in_cim<68>:I 
*.PININFO data_in_cim<67>:I data_in_cim<66>:I data_in_cim<65>:I 
*.PININFO data_in_cim<64>:I data_in_cim<63>:I data_in_cim<62>:I 
*.PININFO data_in_cim<61>:I data_in_cim<60>:I data_in_cim<59>:I 
*.PININFO data_in_cim<58>:I data_in_cim<57>:I data_in_cim<56>:I 
*.PININFO data_in_cim<55>:I data_in_cim<54>:I data_in_cim<53>:I 
*.PININFO data_in_cim<52>:I data_in_cim<51>:I data_in_cim<50>:I 
*.PININFO data_in_cim<49>:I data_in_cim<48>:I data_in_cim<47>:I 
*.PININFO data_in_cim<46>:I data_in_cim<45>:I data_in_cim<44>:I 
*.PININFO data_in_cim<43>:I data_in_cim<42>:I data_in_cim<41>:I 
*.PININFO data_in_cim<40>:I data_in_cim<39>:I data_in_cim<38>:I 
*.PININFO data_in_cim<37>:I data_in_cim<36>:I data_in_cim<35>:I 
*.PININFO data_in_cim<34>:I data_in_cim<33>:I data_in_cim<32>:I 
*.PININFO data_in_cim<31>:I data_in_cim<30>:I data_in_cim<29>:I 
*.PININFO data_in_cim<28>:I data_in_cim<27>:I data_in_cim<26>:I 
*.PININFO data_in_cim<25>:I data_in_cim<24>:I data_in_cim<23>:I 
*.PININFO data_in_cim<22>:I data_in_cim<21>:I data_in_cim<20>:I 
*.PININFO data_in_cim<19>:I data_in_cim<18>:I data_in_cim<17>:I 
*.PININFO data_in_cim<16>:I data_in_cim<15>:I data_in_cim<14>:I 
*.PININFO data_in_cim<13>:I data_in_cim<12>:I data_in_cim<11>:I 
*.PININFO data_in_cim<10>:I data_in_cim<9>:I data_in_cim<8>:I data_in_cim<7>:I 
*.PININFO data_in_cim<6>:I data_in_cim<5>:I data_in_cim<4>:I data_in_cim<3>:I 
*.PININFO data_in_cim<2>:I data_in_cim<1>:I data_in_cim<0>:I inbit:I model:I 
*.PININFO reg_en:I sel_array<15>:I sel_array<14>:I sel_array<13>:I 
*.PININFO sel_array<12>:I sel_array<11>:I sel_array<10>:I sel_array<9>:I 
*.PININFO sel_array<8>:I sel_array<7>:I sel_array<6>:I sel_array<5>:I 
*.PININFO sel_array<4>:I sel_array<3>:I sel_array<2>:I sel_array<1>:I 
*.PININFO sel_array<0>:I set:I wait_:I wrt:I q<191>:O q<190>:O q<189>:O 
*.PININFO q<188>:O q<187>:O q<186>:O q<185>:O q<184>:O q<183>:O q<182>:O 
*.PININFO q<181>:O q<180>:O q<179>:O q<178>:O q<177>:O q<176>:O q<175>:O 
*.PININFO q<174>:O q<173>:O q<172>:O q<171>:O q<170>:O q<169>:O q<168>:O 
*.PININFO q<167>:O q<166>:O q<165>:O q<164>:O q<163>:O q<162>:O q<161>:O 
*.PININFO q<160>:O q<159>:O q<158>:O q<157>:O q<156>:O q<155>:O q<154>:O 
*.PININFO q<153>:O q<152>:O q<151>:O q<150>:O q<149>:O q<148>:O q<147>:O 
*.PININFO q<146>:O q<145>:O q<144>:O q<143>:O q<142>:O q<141>:O q<140>:O 
*.PININFO q<139>:O q<138>:O q<137>:O q<136>:O q<135>:O q<134>:O q<133>:O 
*.PININFO q<132>:O q<131>:O q<130>:O q<129>:O q<128>:O q<127>:O q<126>:O 
*.PININFO q<125>:O q<124>:O q<123>:O q<122>:O q<121>:O q<120>:O q<119>:O 
*.PININFO q<118>:O q<117>:O q<116>:O q<115>:O q<114>:O q<113>:O q<112>:O 
*.PININFO q<111>:O q<110>:O q<109>:O q<108>:O q<107>:O q<106>:O q<105>:O 
*.PININFO q<104>:O q<103>:O q<102>:O q<101>:O q<100>:O q<99>:O q<98>:O q<97>:O 
*.PININFO q<96>:O q<95>:O q<94>:O q<93>:O q<92>:O q<91>:O q<90>:O q<89>:O 
*.PININFO q<88>:O q<87>:O q<86>:O q<85>:O q<84>:O q<83>:O q<82>:O q<81>:O 
*.PININFO q<80>:O q<79>:O q<78>:O q<77>:O q<76>:O q<75>:O q<74>:O q<73>:O 
*.PININFO q<72>:O q<71>:O q<70>:O q<69>:O q<68>:O q<67>:O q<66>:O q<65>:O 
*.PININFO q<64>:O q<63>:O q<62>:O q<61>:O q<60>:O q<59>:O q<58>:O q<57>:O 
*.PININFO q<56>:O q<55>:O q<54>:O q<53>:O q<52>:O q<51>:O q<50>:O q<49>:O 
*.PININFO q<48>:O q<47>:O q<46>:O q<45>:O q<44>:O q<43>:O q<42>:O q<41>:O 
*.PININFO q<40>:O q<39>:O q<38>:O q<37>:O q<36>:O q<35>:O q<34>:O q<33>:O 
*.PININFO q<32>:O q<31>:O q<30>:O q<29>:O q<28>:O q<27>:O q<26>:O q<25>:O 
*.PININFO q<24>:O q<23>:O q<22>:O q<21>:O q<20>:O q<19>:O q<18>:O q<17>:O 
*.PININFO q<16>:O q<15>:O q<14>:O q<13>:O q<12>:O q<11>:O q<10>:O q<9>:O 
*.PININFO q<8>:O q<7>:O q<6>:O q<5>:O q<4>:O q<3>:O q<2>:O q<1>:O q<0>:O vdd:B 
*.PININFO vss:B
XI0 net33<0> net33<1> net33<2> net33<3> net33<4> net33<5> net33<6> net33<7> 
+ net33<8> net33<9> net33<10> net33<11> net33<12> net33<13> net33<14> 
+ net33<15> net33<16> net33<17> net33<18> net33<19> net33<20> net33<21> 
+ net33<22> net33<23> net33<24> net33<25> net33<26> net33<27> net33<28> 
+ net33<29> net33<30> net33<31> net33<32> net33<33> net33<34> net33<35> 
+ net33<36> net33<37> net33<38> net33<39> net33<40> net33<41> net33<42> 
+ net33<43> net33<44> net33<45> net33<46> net33<47> net33<48> net33<49> 
+ net33<50> net33<51> net33<52> net33<53> net33<54> net33<55> net33<56> 
+ net33<57> net33<58> net33<59> net33<60> net33<61> net33<62> net33<63> 
+ net39<0> net39<1> net39<2> net39<3> net39<4> net39<5> net39<6> net39<7> 
+ net39<8> net39<9> net39<10> net39<11> net39<12> net39<13> net39<14> 
+ net39<15> net39<16> net39<17> net39<18> net39<19> net39<20> net39<21> 
+ net39<22> net39<23> net39<24> net39<25> net39<26> net39<27> net39<28> 
+ net39<29> net39<30> net39<31> col_en net31<0> net31<1> net31<2> net31<3> 
+ net31<4> net31<5> net31<6> net31<7> net31<8> net31<9> net31<10> net31<11> 
+ net31<12> net31<13> net31<14> net31<15> net31<16> net31<17> net31<18> 
+ net31<19> net31<20> net31<21> net31<22> net31<23> net31<24> net31<25> 
+ net31<26> net31<27> net31<28> net31<29> net31<30> net31<31> net31<32> 
+ net31<33> net31<34> net31<35> net31<36> net31<37> net31<38> net31<39> 
+ net31<40> net31<41> net31<42> net31<43> net31<44> net31<45> net31<46> 
+ net31<47> net31<48> net31<49> net31<50> net31<51> net31<52> net31<53> 
+ net31<54> net31<55> net31<56> net31<57> net31<58> net31<59> net31<60> 
+ net31<61> net31<62> net31<63> net31<64> net31<65> net31<66> net31<67> 
+ net31<68> net31<69> net31<70> net31<71> net31<72> net31<73> net31<74> 
+ net31<75> net31<76> net31<77> net31<78> net31<79> net31<80> net31<81> 
+ net31<82> net31<83> net31<84> net31<85> net31<86> net31<87> net31<88> 
+ net31<89> net31<90> net31<91> net31<92> net31<93> net31<94> net31<95> 
+ net31<96> net31<97> net31<98> net31<99> net31<100> net31<101> net31<102> 
+ net31<103> net31<104> net31<105> net31<106> net31<107> net31<108> net31<109> 
+ net31<110> net31<111> net31<112> net31<113> net31<114> net31<115> net31<116> 
+ net31<117> net31<118> net31<119> net31<120> net31<121> net31<122> net31<123> 
+ net31<124> net31<125> net31<126> net31<127> net28<0> net28<1> net28<2> 
+ net28<3> net28<4> net28<5> net28<6> net28<7> net28<8> net28<9> net28<10> 
+ net28<11> net28<12> net28<13> net28<14> net28<15> net28<16> net28<17> 
+ net28<18> net28<19> net28<20> net28<21> net28<22> net28<23> net28<24> 
+ net28<25> net28<26> net28<27> net28<28> net28<29> net28<30> net28<31> 
+ net28<32> net28<33> net28<34> net28<35> net28<36> net28<37> net28<38> 
+ net28<39> net28<40> net28<41> net28<42> net28<43> net28<44> net28<45> 
+ net28<46> net28<47> net28<48> net28<49> net28<50> net28<51> net28<52> 
+ net28<53> net28<54> net28<55> net28<56> net28<57> net28<58> net28<59> 
+ net28<60> net28<61> net28<62> net28<63> net28<64> net28<65> net28<66> 
+ net28<67> net28<68> net28<69> net28<70> net28<71> net28<72> net28<73> 
+ net28<74> net28<75> net28<76> net28<77> net28<78> net28<79> net28<80> 
+ net28<81> net28<82> net28<83> net28<84> net28<85> net28<86> net28<87> 
+ net28<88> net28<89> net28<90> net28<91> net28<92> net28<93> net28<94> 
+ net28<95> net28<96> net28<97> net28<98> net28<99> net28<100> net28<101> 
+ net28<102> net28<103> net28<104> net28<105> net28<106> net28<107> net28<108> 
+ net28<109> net28<110> net28<111> net28<112> net28<113> net28<114> net28<115> 
+ net28<116> net28<117> net28<118> net28<119> net28<120> net28<121> net28<122> 
+ net28<123> net28<124> net28<125> net28<126> net28<127> reg_en sel_array<0> 
+ sel_array<1> sel_array<2> sel_array<3> sel_array<4> sel_array<5> 
+ sel_array<6> sel_array<7> sel_array<8> sel_array<9> sel_array<10> 
+ sel_array<11> sel_array<12> sel_array<13> sel_array<14> sel_array<15> 
+ net49<0> net49<1> net49<2> net49<3> net49<4> net49<5> net49<6> net49<7> 
+ net49<8> net49<9> net49<10> net49<11> net49<12> net49<13> net49<14> 
+ net49<15> net49<16> net49<17> net49<18> net49<19> net49<20> net49<21> 
+ net49<22> net49<23> net49<24> net49<25> net49<26> net49<27> net49<28> 
+ net49<29> net49<30> net49<31> net49<32> net49<33> net49<34> net49<35> 
+ net49<36> net49<37> net49<38> net49<39> net49<40> net49<41> net49<42> 
+ net49<43> net49<44> net49<45> net49<46> net49<47> net49<48> net49<49> 
+ net49<50> net49<51> net49<52> net49<53> net49<54> net49<55> net49<56> 
+ net49<57> net49<58> net49<59> net49<60> net49<61> net49<62> net49<63> vdd 
+ vss net35<0> net35<1> net35<2> net35<3> net35<4> net35<5> net35<6> net35<7> 
+ net35<8> net35<9> net35<10> net35<11> net35<12> net35<13> net35<14> 
+ net35<15> net35<16> net35<17> net35<18> net35<19> net35<20> net35<21> 
+ net35<22> net35<23> net35<24> net35<25> net35<26> net35<27> net35<28> 
+ net35<29> net35<30> net35<31> net35<32> net35<33> net35<34> net35<35> 
+ net35<36> net35<37> net35<38> net35<39> net35<40> net35<41> net35<42> 
+ net35<43> net35<44> net35<45> net35<46> net35<47> net35<48> net35<49> 
+ net35<50> net35<51> net35<52> net35<53> net35<54> net35<55> net35<56> 
+ net35<57> net35<58> net35<59> net35<60> net35<61> net35<62> net35<63> 
+ net35<64> net35<65> net35<66> net35<67> net35<68> net35<69> net35<70> 
+ net35<71> net35<72> net35<73> net35<74> net35<75> net35<76> net35<77> 
+ net35<78> net35<79> net35<80> net35<81> net35<82> net35<83> net35<84> 
+ net35<85> net35<86> net35<87> net35<88> net35<89> net35<90> net35<91> 
+ net35<92> net35<93> net35<94> net35<95> net35<96> net35<97> net35<98> 
+ net35<99> net35<100> net35<101> net35<102> net35<103> net35<104> net35<105> 
+ net35<106> net35<107> net35<108> net35<109> net35<110> net35<111> net35<112> 
+ net35<113> net35<114> net35<115> net35<116> net35<117> net35<118> net35<119> 
+ net35<120> net35<121> net35<122> net35<123> net35<124> net35<125> net35<126> 
+ net35<127> / array_test
XI8 net36<0> net36<1> net36<2> net36<3> net36<4> net36<5> net36<6> net36<7> 
+ net36<8> net36<9> net36<10> net36<11> net36<12> net36<13> net36<14> 
+ net36<15> net36<16> net36<17> net36<18> net36<19> net36<20> net36<21> 
+ net36<22> net36<23> net36<24> net36<25> net36<26> net36<27> net36<28> 
+ net36<29> net36<30> net36<31> col_en d<0> d<1> d<2> d<3> d<4> d<5> d<6> d<7> 
+ d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> d<16> d<17> d<18> d<19> d<20> 
+ d<21> d<22> d<23> d<24> d<25> d<26> d<27> d<28> d<29> d<30> d<31> q<0> q<1> 
+ q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> q<15> 
+ q<16> q<17> q<18> q<19> q<20> q<21> q<22> q<23> q<24> q<25> q<26> q<27> 
+ q<28> q<29> q<30> q<31> q<32> q<33> q<34> q<35> q<36> q<37> q<38> q<39> 
+ q<40> q<41> q<42> q<43> q<44> q<45> q<46> q<47> q<48> q<49> q<50> q<51> 
+ q<52> q<53> q<54> q<55> q<56> q<57> q<58> q<59> q<60> q<61> q<62> q<63> 
+ q<64> q<65> q<66> q<67> q<68> q<69> q<70> q<71> q<72> q<73> q<74> q<75> 
+ q<76> q<77> q<78> q<79> q<80> q<81> q<82> q<83> q<84> q<85> q<86> q<87> 
+ q<88> q<89> q<90> q<91> q<92> q<93> q<94> q<95> q<96> q<97> q<98> q<99> 
+ q<100> q<101> q<102> q<103> q<104> q<105> q<106> q<107> q<108> q<109> q<110> 
+ q<111> q<112> q<113> q<114> q<115> q<116> q<117> q<118> q<119> q<120> q<121> 
+ q<122> q<123> q<124> q<125> q<126> q<127> q<128> q<129> q<130> q<131> q<132> 
+ q<133> q<134> q<135> q<136> q<137> q<138> q<139> q<140> q<141> q<142> q<143> 
+ q<144> q<145> q<146> q<147> q<148> q<149> q<150> q<151> q<152> q<153> q<154> 
+ q<155> q<156> q<157> q<158> q<159> q<160> q<161> q<162> q<163> q<164> q<165> 
+ q<166> q<167> q<168> q<169> q<170> q<171> q<172> q<173> q<174> q<175> q<176> 
+ q<177> q<178> q<179> q<180> q<181> q<182> q<183> q<184> q<185> q<186> q<187> 
+ q<188> q<189> q<190> q<191> net41 vdd vss / counter
XI4 a<0> a<1> a<2> a<3> a<4> a<5> a<6> a<7> net46<0> net46<1> net51<0> 
+ net51<1> net51<2> net51<3> net51<4> net51<5> net51<6> clk comp net54 net61 
+ net56 inbit model net40 set net41 net42 net60 net59 net58 net57 vdd vss 
+ wait_ wrt net62 net63 / master
XI11 net36<0> net36<1> net36<2> net36<3> net36<4> net36<5> net36<6> net36<7> 
+ net36<8> net36<9> net36<10> net36<11> net36<12> net36<13> net36<14> 
+ net36<15> net36<16> net36<17> net36<18> net36<19> net36<20> net36<21> 
+ net36<22> net36<23> net36<24> net36<25> net36<26> net36<27> net36<28> 
+ net36<29> net36<30> net36<31> net39<0> net39<1> net39<2> net39<3> net39<4> 
+ net39<5> net39<6> net39<7> net39<8> net39<9> net39<10> net39<11> net39<12> 
+ net39<13> net39<14> net39<15> net39<16> net39<17> net39<18> net39<19> 
+ net39<20> net39<21> net39<22> net39<23> net39<24> net39<25> net39<26> 
+ net39<27> net39<28> net39<29> net39<30> net39<31> d<0> d<1> d<2> d<3> d<4> 
+ d<5> d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> d<16> d<17> 
+ d<18> d<19> d<20> d<21> d<22> d<23> d<24> d<25> d<26> d<27> d<28> d<29> 
+ d<30> d<31> net40 net41 net42 vdd vss / ADC
XI2 net33<0> net33<1> net33<2> net33<3> net33<4> net33<5> net33<6> net33<7> 
+ net33<8> net33<9> net33<10> net33<11> net33<12> net33<13> net33<14> 
+ net33<15> net33<16> net33<17> net33<18> net33<19> net33<20> net33<21> 
+ net33<22> net33<23> net33<24> net33<25> net33<26> net33<27> net33<28> 
+ net33<29> net33<30> net33<31> net33<32> net33<33> net33<34> net33<35> 
+ net33<36> net33<37> net33<38> net33<39> net33<40> net33<41> net33<42> 
+ net33<43> net33<44> net33<45> net33<46> net33<47> net33<48> net33<49> 
+ net33<50> net33<51> net33<52> net33<53> net33<54> net33<55> net33<56> 
+ net33<57> net33<58> net33<59> net33<60> net33<61> net33<62> net33<63> 
+ net39<0> net39<1> net39<2> net39<3> net39<4> net39<5> net39<6> net39<7> 
+ net39<8> net39<9> net39<10> net39<11> net39<12> net39<13> net39<14> 
+ net39<15> net39<16> net39<17> net39<18> net39<19> net39<20> net39<21> 
+ net39<22> net39<23> net39<24> net39<25> net39<26> net39<27> net39<28> 
+ net39<29> net39<30> net39<31> net012<0> net012<1> d<0> d<1> d<2> d<3> d<4> 
+ d<5> d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> d<16> d<17> 
+ d<18> d<19> d<20> d<21> d<22> d<23> d<24> d<25> d<26> d<27> d<28> d<29> 
+ d<30> d<31> reg_en net49<0> net49<1> net49<2> net49<3> net49<4> net49<5> 
+ net49<6> net49<7> net49<8> net49<9> net49<10> net49<11> net49<12> net49<13> 
+ net49<14> net49<15> net49<16> net49<17> net49<18> net49<19> net49<20> 
+ net49<21> net49<22> net49<23> net49<24> net49<25> net49<26> net49<27> 
+ net49<28> net49<29> net49<30> net49<31> net49<32> net49<33> net49<34> 
+ net49<35> net49<36> net49<37> net49<38> net49<39> net49<40> net49<41> 
+ net49<42> net49<43> net49<44> net49<45> net49<46> net49<47> net49<48> 
+ net49<49> net49<50> net49<51> net49<52> net49<53> net49<54> net49<55> 
+ net49<56> net49<57> net49<58> net49<59> net49<60> net49<61> net49<62> 
+ net49<63> vdd vss net62 net63 / Writedriver
XI3 net46<0> net46<1> net51<0> net51<1> net51<2> net51<3> net51<4> net51<5> 
+ net51<6> net012<0> net012<1> net54 net61 net45<0> net45<1> net45<2> net45<3> 
+ net45<4> net45<5> net45<6> net45<7> reg_en net44<0> net44<1> net44<2> 
+ net44<3> net44<4> net44<5> net44<6> net44<7> net44<8> net44<9> net44<10> 
+ net44<11> net44<12> net44<13> net44<14> net44<15> vdd vss net62 net63 / 
+ access_decoder
XI7 net56 net31<0> net31<1> net31<2> net31<3> net31<4> net31<5> net31<6> 
+ net31<7> net31<8> net31<9> net31<10> net31<11> net31<12> net31<13> net31<14> 
+ net31<15> net31<16> net31<17> net31<18> net31<19> net31<20> net31<21> 
+ net31<22> net31<23> net31<24> net31<25> net31<26> net31<27> net31<28> 
+ net31<29> net31<30> net31<31> net31<32> net31<33> net31<34> net31<35> 
+ net31<36> net31<37> net31<38> net31<39> net31<40> net31<41> net31<42> 
+ net31<43> net31<44> net31<45> net31<46> net31<47> net31<48> net31<49> 
+ net31<50> net31<51> net31<52> net31<53> net31<54> net31<55> net31<56> 
+ net31<57> net31<58> net31<59> net31<60> net31<61> net31<62> net31<63> 
+ net31<64> net31<65> net31<66> net31<67> net31<68> net31<69> net31<70> 
+ net31<71> net31<72> net31<73> net31<74> net31<75> net31<76> net31<77> 
+ net31<78> net31<79> net31<80> net31<81> net31<82> net31<83> net31<84> 
+ net31<85> net31<86> net31<87> net31<88> net31<89> net31<90> net31<91> 
+ net31<92> net31<93> net31<94> net31<95> net31<96> net31<97> net31<98> 
+ net31<99> net31<100> net31<101> net31<102> net31<103> net31<104> net31<105> 
+ net31<106> net31<107> net31<108> net31<109> net31<110> net31<111> net31<112> 
+ net31<113> net31<114> net31<115> net31<116> net31<117> net31<118> net31<119> 
+ net31<120> net31<121> net31<122> net31<123> net31<124> net31<125> net31<126> 
+ net31<127> net28<0> net28<1> net28<2> net28<3> net28<4> net28<5> net28<6> 
+ net28<7> net28<8> net28<9> net28<10> net28<11> net28<12> net28<13> net28<14> 
+ net28<15> net28<16> net28<17> net28<18> net28<19> net28<20> net28<21> 
+ net28<22> net28<23> net28<24> net28<25> net28<26> net28<27> net28<28> 
+ net28<29> net28<30> net28<31> net28<32> net28<33> net28<34> net28<35> 
+ net28<36> net28<37> net28<38> net28<39> net28<40> net28<41> net28<42> 
+ net28<43> net28<44> net28<45> net28<46> net28<47> net28<48> net28<49> 
+ net28<50> net28<51> net28<52> net28<53> net28<54> net28<55> net28<56> 
+ net28<57> net28<58> net28<59> net28<60> net28<61> net28<62> net28<63> 
+ net28<64> net28<65> net28<66> net28<67> net28<68> net28<69> net28<70> 
+ net28<71> net28<72> net28<73> net28<74> net28<75> net28<76> net28<77> 
+ net28<78> net28<79> net28<80> net28<81> net28<82> net28<83> net28<84> 
+ net28<85> net28<86> net28<87> net28<88> net28<89> net28<90> net28<91> 
+ net28<92> net28<93> net28<94> net28<95> net28<96> net28<97> net28<98> 
+ net28<99> net28<100> net28<101> net28<102> net28<103> net28<104> net28<105> 
+ net28<106> net28<107> net28<108> net28<109> net28<110> net28<111> net28<112> 
+ net28<113> net28<114> net28<115> net28<116> net28<117> net28<118> net28<119> 
+ net28<120> net28<121> net28<122> net28<123> net28<124> net28<125> net28<126> 
+ net28<127> data_in_cim<0> data_in_cim<1> data_in_cim<2> data_in_cim<3> 
+ data_in_cim<4> data_in_cim<5> data_in_cim<6> data_in_cim<7> data_in_cim<8> 
+ data_in_cim<9> data_in_cim<10> data_in_cim<11> data_in_cim<12> 
+ data_in_cim<13> data_in_cim<14> data_in_cim<15> data_in_cim<16> 
+ data_in_cim<17> data_in_cim<18> data_in_cim<19> data_in_cim<20> 
+ data_in_cim<21> data_in_cim<22> data_in_cim<23> data_in_cim<24> 
+ data_in_cim<25> data_in_cim<26> data_in_cim<27> data_in_cim<28> 
+ data_in_cim<29> data_in_cim<30> data_in_cim<31> data_in_cim<32> 
+ data_in_cim<33> data_in_cim<34> data_in_cim<35> data_in_cim<36> 
+ data_in_cim<37> data_in_cim<38> data_in_cim<39> data_in_cim<40> 
+ data_in_cim<41> data_in_cim<42> data_in_cim<43> data_in_cim<44> 
+ data_in_cim<45> data_in_cim<46> data_in_cim<47> data_in_cim<48> 
+ data_in_cim<49> data_in_cim<50> data_in_cim<51> data_in_cim<52> 
+ data_in_cim<53> data_in_cim<54> data_in_cim<55> data_in_cim<56> 
+ data_in_cim<57> data_in_cim<58> data_in_cim<59> data_in_cim<60> 
+ data_in_cim<61> data_in_cim<62> data_in_cim<63> data_in_cim<64> 
+ data_in_cim<65> data_in_cim<66> data_in_cim<67> data_in_cim<68> 
+ data_in_cim<69> data_in_cim<70> data_in_cim<71> data_in_cim<72> 
+ data_in_cim<73> data_in_cim<74> data_in_cim<75> data_in_cim<76> 
+ data_in_cim<77> data_in_cim<78> data_in_cim<79> data_in_cim<80> 
+ data_in_cim<81> data_in_cim<82> data_in_cim<83> data_in_cim<84> 
+ data_in_cim<85> data_in_cim<86> data_in_cim<87> data_in_cim<88> 
+ data_in_cim<89> data_in_cim<90> data_in_cim<91> data_in_cim<92> 
+ data_in_cim<93> data_in_cim<94> data_in_cim<95> data_in_cim<96> 
+ data_in_cim<97> data_in_cim<98> data_in_cim<99> data_in_cim<100> 
+ data_in_cim<101> data_in_cim<102> data_in_cim<103> data_in_cim<104> 
+ data_in_cim<105> data_in_cim<106> data_in_cim<107> data_in_cim<108> 
+ data_in_cim<109> data_in_cim<110> data_in_cim<111> data_in_cim<112> 
+ data_in_cim<113> data_in_cim<114> data_in_cim<115> data_in_cim<116> 
+ data_in_cim<117> data_in_cim<118> data_in_cim<119> data_in_cim<120> 
+ data_in_cim<121> data_in_cim<122> data_in_cim<123> data_in_cim<124> 
+ data_in_cim<125> data_in_cim<126> data_in_cim<127> data_in_cim<128> 
+ data_in_cim<129> data_in_cim<130> data_in_cim<131> data_in_cim<132> 
+ data_in_cim<133> data_in_cim<134> data_in_cim<135> data_in_cim<136> 
+ data_in_cim<137> data_in_cim<138> data_in_cim<139> data_in_cim<140> 
+ data_in_cim<141> data_in_cim<142> data_in_cim<143> data_in_cim<144> 
+ data_in_cim<145> data_in_cim<146> data_in_cim<147> data_in_cim<148> 
+ data_in_cim<149> data_in_cim<150> data_in_cim<151> data_in_cim<152> 
+ data_in_cim<153> data_in_cim<154> data_in_cim<155> data_in_cim<156> 
+ data_in_cim<157> data_in_cim<158> data_in_cim<159> data_in_cim<160> 
+ data_in_cim<161> data_in_cim<162> data_in_cim<163> data_in_cim<164> 
+ data_in_cim<165> data_in_cim<166> data_in_cim<167> data_in_cim<168> 
+ data_in_cim<169> data_in_cim<170> data_in_cim<171> data_in_cim<172> 
+ data_in_cim<173> data_in_cim<174> data_in_cim<175> data_in_cim<176> 
+ data_in_cim<177> data_in_cim<178> data_in_cim<179> data_in_cim<180> 
+ data_in_cim<181> data_in_cim<182> data_in_cim<183> data_in_cim<184> 
+ data_in_cim<185> data_in_cim<186> data_in_cim<187> data_in_cim<188> 
+ data_in_cim<189> data_in_cim<190> data_in_cim<191> data_in_cim<192> 
+ data_in_cim<193> data_in_cim<194> data_in_cim<195> data_in_cim<196> 
+ data_in_cim<197> data_in_cim<198> data_in_cim<199> data_in_cim<200> 
+ data_in_cim<201> data_in_cim<202> data_in_cim<203> data_in_cim<204> 
+ data_in_cim<205> data_in_cim<206> data_in_cim<207> data_in_cim<208> 
+ data_in_cim<209> data_in_cim<210> data_in_cim<211> data_in_cim<212> 
+ data_in_cim<213> data_in_cim<214> data_in_cim<215> data_in_cim<216> 
+ data_in_cim<217> data_in_cim<218> data_in_cim<219> data_in_cim<220> 
+ data_in_cim<221> data_in_cim<222> data_in_cim<223> data_in_cim<224> 
+ data_in_cim<225> data_in_cim<226> data_in_cim<227> data_in_cim<228> 
+ data_in_cim<229> data_in_cim<230> data_in_cim<231> data_in_cim<232> 
+ data_in_cim<233> data_in_cim<234> data_in_cim<235> data_in_cim<236> 
+ data_in_cim<237> data_in_cim<238> data_in_cim<239> data_in_cim<240> 
+ data_in_cim<241> data_in_cim<242> data_in_cim<243> data_in_cim<244> 
+ data_in_cim<245> data_in_cim<246> data_in_cim<247> data_in_cim<248> 
+ data_in_cim<249> data_in_cim<250> data_in_cim<251> data_in_cim<252> 
+ data_in_cim<253> data_in_cim<254> data_in_cim<255> data_in_cim<256> 
+ data_in_cim<257> data_in_cim<258> data_in_cim<259> data_in_cim<260> 
+ data_in_cim<261> data_in_cim<262> data_in_cim<263> data_in_cim<264> 
+ data_in_cim<265> data_in_cim<266> data_in_cim<267> data_in_cim<268> 
+ data_in_cim<269> data_in_cim<270> data_in_cim<271> data_in_cim<272> 
+ data_in_cim<273> data_in_cim<274> data_in_cim<275> data_in_cim<276> 
+ data_in_cim<277> data_in_cim<278> data_in_cim<279> data_in_cim<280> 
+ data_in_cim<281> data_in_cim<282> data_in_cim<283> data_in_cim<284> 
+ data_in_cim<285> data_in_cim<286> data_in_cim<287> data_in_cim<288> 
+ data_in_cim<289> data_in_cim<290> data_in_cim<291> data_in_cim<292> 
+ data_in_cim<293> data_in_cim<294> data_in_cim<295> data_in_cim<296> 
+ data_in_cim<297> data_in_cim<298> data_in_cim<299> data_in_cim<300> 
+ data_in_cim<301> data_in_cim<302> data_in_cim<303> data_in_cim<304> 
+ data_in_cim<305> data_in_cim<306> data_in_cim<307> data_in_cim<308> 
+ data_in_cim<309> data_in_cim<310> data_in_cim<311> data_in_cim<312> 
+ data_in_cim<313> data_in_cim<314> data_in_cim<315> data_in_cim<316> 
+ data_in_cim<317> data_in_cim<318> data_in_cim<319> data_in_cim<320> 
+ data_in_cim<321> data_in_cim<322> data_in_cim<323> data_in_cim<324> 
+ data_in_cim<325> data_in_cim<326> data_in_cim<327> data_in_cim<328> 
+ data_in_cim<329> data_in_cim<330> data_in_cim<331> data_in_cim<332> 
+ data_in_cim<333> data_in_cim<334> data_in_cim<335> data_in_cim<336> 
+ data_in_cim<337> data_in_cim<338> data_in_cim<339> data_in_cim<340> 
+ data_in_cim<341> data_in_cim<342> data_in_cim<343> data_in_cim<344> 
+ data_in_cim<345> data_in_cim<346> data_in_cim<347> data_in_cim<348> 
+ data_in_cim<349> data_in_cim<350> data_in_cim<351> data_in_cim<352> 
+ data_in_cim<353> data_in_cim<354> data_in_cim<355> data_in_cim<356> 
+ data_in_cim<357> data_in_cim<358> data_in_cim<359> data_in_cim<360> 
+ data_in_cim<361> data_in_cim<362> data_in_cim<363> data_in_cim<364> 
+ data_in_cim<365> data_in_cim<366> data_in_cim<367> data_in_cim<368> 
+ data_in_cim<369> data_in_cim<370> data_in_cim<371> data_in_cim<372> 
+ data_in_cim<373> data_in_cim<374> data_in_cim<375> data_in_cim<376> 
+ data_in_cim<377> data_in_cim<378> data_in_cim<379> data_in_cim<380> 
+ data_in_cim<381> data_in_cim<382> data_in_cim<383> data_in_cim<384> 
+ data_in_cim<385> data_in_cim<386> data_in_cim<387> data_in_cim<388> 
+ data_in_cim<389> data_in_cim<390> data_in_cim<391> data_in_cim<392> 
+ data_in_cim<393> data_in_cim<394> data_in_cim<395> data_in_cim<396> 
+ data_in_cim<397> data_in_cim<398> data_in_cim<399> data_in_cim<400> 
+ data_in_cim<401> data_in_cim<402> data_in_cim<403> data_in_cim<404> 
+ data_in_cim<405> data_in_cim<406> data_in_cim<407> data_in_cim<408> 
+ data_in_cim<409> data_in_cim<410> data_in_cim<411> data_in_cim<412> 
+ data_in_cim<413> data_in_cim<414> data_in_cim<415> data_in_cim<416> 
+ data_in_cim<417> data_in_cim<418> data_in_cim<419> data_in_cim<420> 
+ data_in_cim<421> data_in_cim<422> data_in_cim<423> data_in_cim<424> 
+ data_in_cim<425> data_in_cim<426> data_in_cim<427> data_in_cim<428> 
+ data_in_cim<429> data_in_cim<430> data_in_cim<431> data_in_cim<432> 
+ data_in_cim<433> data_in_cim<434> data_in_cim<435> data_in_cim<436> 
+ data_in_cim<437> data_in_cim<438> data_in_cim<439> data_in_cim<440> 
+ data_in_cim<441> data_in_cim<442> data_in_cim<443> data_in_cim<444> 
+ data_in_cim<445> data_in_cim<446> data_in_cim<447> data_in_cim<448> 
+ data_in_cim<449> data_in_cim<450> data_in_cim<451> data_in_cim<452> 
+ data_in_cim<453> data_in_cim<454> data_in_cim<455> data_in_cim<456> 
+ data_in_cim<457> data_in_cim<458> data_in_cim<459> data_in_cim<460> 
+ data_in_cim<461> data_in_cim<462> data_in_cim<463> data_in_cim<464> 
+ data_in_cim<465> data_in_cim<466> data_in_cim<467> data_in_cim<468> 
+ data_in_cim<469> data_in_cim<470> data_in_cim<471> data_in_cim<472> 
+ data_in_cim<473> data_in_cim<474> data_in_cim<475> data_in_cim<476> 
+ data_in_cim<477> data_in_cim<478> data_in_cim<479> data_in_cim<480> 
+ data_in_cim<481> data_in_cim<482> data_in_cim<483> data_in_cim<484> 
+ data_in_cim<485> data_in_cim<486> data_in_cim<487> data_in_cim<488> 
+ data_in_cim<489> data_in_cim<490> data_in_cim<491> data_in_cim<492> 
+ data_in_cim<493> data_in_cim<494> data_in_cim<495> data_in_cim<496> 
+ data_in_cim<497> data_in_cim<498> data_in_cim<499> data_in_cim<500> 
+ data_in_cim<501> data_in_cim<502> data_in_cim<503> data_in_cim<504> 
+ data_in_cim<505> data_in_cim<506> data_in_cim<507> data_in_cim<508> 
+ data_in_cim<509> data_in_cim<510> data_in_cim<511> net60 net59 net58 net57 
+ vdd vss / timegenerate
XI10 net45<0> net45<1> net45<2> net45<3> net45<4> net45<5> net45<6> net45<7> 
+ net31<0> net31<1> net31<2> net31<3> net31<4> net31<5> net31<6> net31<7> 
+ net31<8> net31<9> net31<10> net31<11> net31<12> net31<13> net31<14> 
+ net31<15> net31<16> net31<17> net31<18> net31<19> net31<20> net31<21> 
+ net31<22> net31<23> net31<24> net31<25> net31<26> net31<27> net31<28> 
+ net31<29> net31<30> net31<31> net31<32> net31<33> net31<34> net31<35> 
+ net31<36> net31<37> net31<38> net31<39> net31<40> net31<41> net31<42> 
+ net31<43> net31<44> net31<45> net31<46> net31<47> net31<48> net31<49> 
+ net31<50> net31<51> net31<52> net31<53> net31<54> net31<55> net31<56> 
+ net31<57> net31<58> net31<59> net31<60> net31<61> net31<62> net31<63> 
+ net31<64> net31<65> net31<66> net31<67> net31<68> net31<69> net31<70> 
+ net31<71> net31<72> net31<73> net31<74> net31<75> net31<76> net31<77> 
+ net31<78> net31<79> net31<80> net31<81> net31<82> net31<83> net31<84> 
+ net31<85> net31<86> net31<87> net31<88> net31<89> net31<90> net31<91> 
+ net31<92> net31<93> net31<94> net31<95> net31<96> net31<97> net31<98> 
+ net31<99> net31<100> net31<101> net31<102> net31<103> net31<104> net31<105> 
+ net31<106> net31<107> net31<108> net31<109> net31<110> net31<111> net31<112> 
+ net31<113> net31<114> net31<115> net31<116> net31<117> net31<118> net31<119> 
+ net31<120> net31<121> net31<122> net31<123> net31<124> net31<125> net31<126> 
+ net31<127> net28<0> net28<1> net28<2> net28<3> net28<4> net28<5> net28<6> 
+ net28<7> net28<8> net28<9> net28<10> net28<11> net28<12> net28<13> net28<14> 
+ net28<15> net28<16> net28<17> net28<18> net28<19> net28<20> net28<21> 
+ net28<22> net28<23> net28<24> net28<25> net28<26> net28<27> net28<28> 
+ net28<29> net28<30> net28<31> net28<32> net28<33> net28<34> net28<35> 
+ net28<36> net28<37> net28<38> net28<39> net28<40> net28<41> net28<42> 
+ net28<43> net28<44> net28<45> net28<46> net28<47> net28<48> net28<49> 
+ net28<50> net28<51> net28<52> net28<53> net28<54> net28<55> net28<56> 
+ net28<57> net28<58> net28<59> net28<60> net28<61> net28<62> net28<63> 
+ net28<64> net28<65> net28<66> net28<67> net28<68> net28<69> net28<70> 
+ net28<71> net28<72> net28<73> net28<74> net28<75> net28<76> net28<77> 
+ net28<78> net28<79> net28<80> net28<81> net28<82> net28<83> net28<84> 
+ net28<85> net28<86> net28<87> net28<88> net28<89> net28<90> net28<91> 
+ net28<92> net28<93> net28<94> net28<95> net28<96> net28<97> net28<98> 
+ net28<99> net28<100> net28<101> net28<102> net28<103> net28<104> net28<105> 
+ net28<106> net28<107> net28<108> net28<109> net28<110> net28<111> net28<112> 
+ net28<113> net28<114> net28<115> net28<116> net28<117> net28<118> net28<119> 
+ net28<120> net28<121> net28<122> net28<123> net28<124> net28<125> net28<126> 
+ net28<127> net44<0> net44<1> net44<2> net44<3> net44<4> net44<5> net44<6> 
+ net44<7> net44<8> net44<9> net44<10> net44<11> net44<12> net44<13> net44<14> 
+ net44<15> vdd vss net35<0> net35<1> net35<2> net35<3> net35<4> net35<5> 
+ net35<6> net35<7> net35<8> net35<9> net35<10> net35<11> net35<12> net35<13> 
+ net35<14> net35<15> net35<16> net35<17> net35<18> net35<19> net35<20> 
+ net35<21> net35<22> net35<23> net35<24> net35<25> net35<26> net35<27> 
+ net35<28> net35<29> net35<30> net35<31> net35<32> net35<33> net35<34> 
+ net35<35> net35<36> net35<37> net35<38> net35<39> net35<40> net35<41> 
+ net35<42> net35<43> net35<44> net35<45> net35<46> net35<47> net35<48> 
+ net35<49> net35<50> net35<51> net35<52> net35<53> net35<54> net35<55> 
+ net35<56> net35<57> net35<58> net35<59> net35<60> net35<61> net35<62> 
+ net35<63> net35<64> net35<65> net35<66> net35<67> net35<68> net35<69> 
+ net35<70> net35<71> net35<72> net35<73> net35<74> net35<75> net35<76> 
+ net35<77> net35<78> net35<79> net35<80> net35<81> net35<82> net35<83> 
+ net35<84> net35<85> net35<86> net35<87> net35<88> net35<89> net35<90> 
+ net35<91> net35<92> net35<93> net35<94> net35<95> net35<96> net35<97> 
+ net35<98> net35<99> net35<100> net35<101> net35<102> net35<103> net35<104> 
+ net35<105> net35<106> net35<107> net35<108> net35<109> net35<110> net35<111> 
+ net35<112> net35<113> net35<114> net35<115> net35<116> net35<117> net35<118> 
+ net35<119> net35<120> net35<121> net35<122> net35<123> net35<124> net35<125> 
+ net35<126> net35<127> / WLdriver_editable

.global vdd vss
v_vss vss 0 0
vsu vdd vss 1.2
*.print v(*)

.ENDS

