* 
* No part of this file can be released without the consent of SMIC.
*
************************************************************************************************************
* smic 0.18um mixed signal 1p6m 1.8v/3.3v spice model(for HSPICE only) *
************************************************************************************************************
*
* Release version    : 1.11
*
* Release date       : 19/03/2015
*
* Simulation tool    : Synopsys Star-HSPICE version C-2009.09
*
*  Inductor   :
* *  *------------------------*---------------------------------------------------------*
*    |  Turn, Radius & Width  |  T=2~7.5 step 0.5,W=3~15um,R=1.7071*W+11.878~120um       |
* *  *------------------------*---------------------------------------------------------*
*    |        Model Name      |              diff_ind_3t_rf_psub                           |
* *  *------------------------*---------------------------------------------------------*
.subckt diff_ind_3t_rf_psub PLUS MINUS CT PSUB R=6e-05 w=8e-06 n=3
.param radius_='0.00833333*(R/1e-06-0)' w_='0.0666667*(w/1e-06-0)'
.param T54='(1-abs(sgn(n-(2.5))))'
.param T55='(min(sgn(radius_-(0.416958))+1,1))'
.param T56='(min(sgn(w_-(0.6004))+1,1))'
.param T57='(min(sgn(w_-(0.5996))+1,1))'
.param T58='(min(sgn(radius_-(0.416375))+1,1))'
.param T59='(min(sgn(radius_-(0.708625))+1,1))'
.param T60='(min(sgn(radius_-(0.708042))+1,1))'
.param T61='(1-abs(sgn(n-(2))))'
.param T62='(1-abs(sgn(n-(3.5))))'
.param T63='(1-abs(sgn(n-(3))))'
.param T64='(1-abs(sgn(n-(4.5))))'
.param T65='(1-abs(sgn(n-(4))))'
.param T66='(1-abs(sgn(n-(5.5))))'
.param T67='(1-abs(sgn(n-(5))))'
.param T68='(1-abs(sgn(n-(6.5))))'
.param T69='(1-abs(sgn(n-(6))))'
.param T70='(1-abs(sgn(n-(7.5))))'
.param T71='(1-abs(sgn(n-(7))))'
.param S0='T54*(1-T55)*(1-T56)'
.param noS0='(1-S0)'
.param S1='T54*T57*(1-T55)*noS0'
.param noS1='(1-S1)*noS0'
.param S2='T54*(1-T56)*T58*(1-T59)*noS1'
.param noS2='(1-S2)*noS1'
.param S3='T54*T58*T57*(1-T59)*noS2'
.param noS3='(1-S3)*noS2'
.param S4='T54*(1-T56)*T60*noS3'
.param noS4='(1-S4)*noS3'
.param S5='T54*T60*T57*noS4'
.param noS5='(1-S5)*noS4'
.param S6='T61*(1-T55)*(1-T56)*noS5'
.param noS6='(1-S6)*noS5'
.param S7='T61*T57*(1-T55)*noS6'
.param noS7='(1-S7)*noS6'
.param S8='T61*(1-T56)*T58*(1-T59)*noS7'
.param noS8='(1-S8)*noS7'
.param S9='T61*T58*T57*(1-T59)*noS8'
.param noS9='(1-S9)*noS8'
.param S10='T61*(1-T56)*T60*noS9'
.param noS10='(1-S10)*noS9'
.param S11='T61*T60*T57*noS10'
.param noS11='(1-S11)*noS10'
.param S12='T62*(1-T55)*noS11'
.param noS12='(1-S12)*noS11'
.param S13='T62*T58*(1-T59)*noS12'
.param noS13='(1-S13)*noS12'
.param S14='T62*T60*noS13'
.param noS14='(1-S14)*noS13'
.param S15='T63*(1-T55)*(1-T56)*noS14'
.param noS15='(1-S15)*noS14'
.param S16='T63*T57*(1-T55)*noS15'
.param noS16='(1-S16)*noS15'
.param S17='T63*(1-T56)*T58*(1-T59)*noS16'
.param noS17='(1-S17)*noS16'
.param S18='T63*T58*T57*(1-T59)*noS17'
.param noS18='(1-S18)*noS17'
.param S19='T63*(1-T56)*T60*noS18'
.param noS19='(1-S19)*noS18'
.param S20='T63*T60*T57*noS19'
.param noS20='(1-S20)*noS19'
.param S21='T64*(1-T55)*noS20'
.param noS21='(1-S21)*noS20'
.param S22='T64*T58*(1-T59)*noS21'
.param noS22='(1-S22)*noS21'
.param S23='T64*T60*noS22'
.param noS23='(1-S23)*noS22'
.param S24='T65*(1-T55)*noS23'
.param noS24='(1-S24)*noS23'
.param S25='T65*T58*(1-T59)*noS24'
.param noS25='(1-S25)*noS24'
.param S26='T65*T60*noS25'
.param noS26='(1-S26)*noS25'
.param S27='T66*(1-T55)*noS26'
.param noS27='(1-S27)*noS26'
.param S28='T66*T58*(1-T59)*noS27'
.param noS28='(1-S28)*noS27'
.param S29='T66*T60*noS28'
.param noS29='(1-S29)*noS28'
.param S30='T67*(1-T55)*noS29'
.param noS30='(1-S30)*noS29'
.param S31='T67*T58*(1-T59)*noS30'
.param noS31='(1-S31)*noS30'
.param S32='T67*T60*noS31'
.param noS32='(1-S32)*noS31'
.param S33='T68*(1-T55)*noS32'
.param noS33='(1-S33)*noS32'
.param S34='T68*T58*(1-T59)*noS33'
.param noS34='(1-S34)*noS33'
.param S35='T68*T60*noS34'
.param noS35='(1-S35)*noS34'
.param S36='T69*(1-T55)*noS35'
.param noS36='(1-S36)*noS35'
.param S37='T69*T58*(1-T59)*noS36'
.param noS37='(1-S37)*noS36'
.param S38='T69*T60*noS37'
.param noS38='(1-S38)*noS37'
.param S39='T70*(1-T55)*noS38'
.param noS39='(1-S39)*noS38'
.param S40='T70*T58*(1-T59)*noS39'
.param noS40='(1-S40)*noS39'
.param S41='T70*T60*noS40'
.param noS41='(1-S41)*noS40'
.param S42='T71*(1-T55)*noS41'
.param noS42='(1-S42)*noS41'
.param S43='T71*T58*(1-T59)*noS42'
.param noS43='(1-S43)*noS42'
.param S44='T71*T60*noS43'
.param noS44='(1-S44)*noS43'
.param V0_part1='7.252626e-03*S0+9.835335e-04*S1+(-9.872708e+00)*S2+5.926542e+00*S3+1.018879e-01*S4+(-8.510330e-03)*S5+(-1.385541e-02)*S6+4.825201e+00*S7+7.062424e-03*S8+1.250880e-01*S9'
.param V0_part2='V0_part1+(-1.097562e-02)*S10+1.035813e-02*S11+(-1.361625e-02)*S12+6.094989e-02*S13+8.011102e-02*S14+2.366697e-01*S15+(-2.694565e-02)*S16+1.519671e+01*S17+5.902280e+00*S18+9.199964e-02*S19'
.param V0_part3='V0_part2+(-6.656587e-03)*S20+4.678773e-02*S21+(-9.423988e+01)*S22+1.380206e+00*S23+(-9.922798e+00)*S24+(-2.388826e+01)*S25+6.909048e-01*S26+(-1.802162e+01)*S27+(-4.314605e+00)*S28+(-1.039441e+01)*S29'
.param V0_part4='V0_part3+(-8.476416e+00)*S30+(-6.694727e+00)*S31+(-3.645804e+00)*S32+(-1.252296e+01)*S33+(-1.415597e+00)*S34+2.758558e+00*S35+(-9.408545e-01)*S36+(-3.027198e+00)*S37+(-1.068115e+01)*S38+(-7.134941e-01)*S39'
.param V0='V0_part4+4.333709e-01*S40+(-1.164668e+01)*S41+8.410414e-01*S42+(-5.467395e+00)*S43+(-1.117661e+01)*S44'
.param V1_part1='9.287330e-01*S0+9.441311e-01*S1+4.210706e+01*S2+3.743246e+01*S3+1.161998e+00*S4+1.116103e+00*S5+6.394954e-01*S6+7.453498e+01*S7+6.513820e-01*S8+2.704156e+01*S9'
.param V1_part2='V1_part1+7.352763e-01*S10+6.476564e-01*S11+1.757831e+00*S12+1.903521e+00*S13+2.088816e+00*S14+4.541104e+01*S15+1.079917e+00*S16+5.007497e+01*S17+3.058275e+01*S18+1.517219e+00*S19'
.param V1_part3='V1_part2+1.430437e+00*S20+2.619119e+00*S21+2.399574e+02*S22+3.168481e+00*S23+2.656848e+02*S24+7.207280e+01*S25+2.883046e+00*S26+1.906885e+02*S27+1.813902e+01*S28+2.820510e+01*S29'
.param V1_part4='V1_part3+1.130780e+02*S30+2.507566e+01*S31+1.233099e+01*S32+2.347975e+02*S33+1.016453e+01*S34+5.812620e+00*S35+1.080422e+01*S36+1.416689e+01*S37+2.734311e+01*S38+1.415998e+01*S39'
.param V1='V1_part4+7.075231e+00*S40+2.939331e+01*S41+9.233226e+00*S42+2.480002e+01*S43+3.116811e+01*S44'
.param V2_part1='(-3.545067e-02)*S0+1.220135e-02*S1+7.265747e-01*S2+(-1.263018e+01)*S3+(-3.304903e-01)*S4+(-1.044161e-01)*S5+(-2.357017e-02)*S6+(-4.836521e+00)*S7+(-7.686143e-02)*S8+(-4.046034e+00)*S9'
.param V2_part2='V2_part1+(-1.506826e-01)*S10+(-8.883717e-02)*S11+3.689071e-02*S12+(-2.584577e-01)*S13+(-5.457140e-01)*S14+(-1.057582e+01)*S15+1.048975e-02*S16+(-2.183820e+01)*S17+(-1.204339e+01)*S18+(-3.841456e-01)*S19'
.param V2_part3='V2_part2+(-1.073917e-01)*S20+1.360732e-02*S21+1.231204e+02*S22+(-1.224182e+00)*S23+(-6.428356e+01)*S24+2.473023e+01*S25+(-1.652991e+00)*S26+6.684535e+00*S27+5.365296e+00*S28+1.115884e+00*S29'
.param V2_part4='V2_part3+(-8.260474e+00)*S30+1.112139e+01*S31+(-3.634629e-01)*S32+(-2.561237e+01)*S33+1.640519e+00*S34+(-2.567087e+00)*S35+3.629807e+00*S36+4.183097e+00*S37+2.639454e+00*S38+2.212107e+00*S39'
.param V2='V2_part4+(-5.010167e-01)*S40+9.821027e+00*S41+(-6.556497e-01)*S42+7.107068e+00*S43+3.401330e-01*S44'
.param V3_part1='(-4.055604e-01)*S0+(-2.154492e-01)*S1+(-1.480783e+02)*S2+(-4.453605e+02)*S3+(-1.484691e+00)*S4+(-7.412859e-01)*S5+(-3.305775e-01)*S6+(-4.536123e+01)*S7+(-6.287504e-01)*S8+(-1.610935e+01)*S9'
.param V3_part2='V3_part1+(-1.059010e+00)*S10+(-5.896743e-01)*S11+(-5.427298e-01)*S12+(-1.404503e+00)*S13+(-2.270820e+00)*S14+(-5.454435e+02)*S15+(-1.929044e-01)*S16+(-9.471442e+01)*S17+(-2.024725e+02)*S18+(-1.677399e+00)*S19'
.param V3_part3='V3_part2+(-8.322557e-01)*S20+(-5.107707e-01)*S21+3.269585e+02*S22+(-3.711010e+00)*S23+(-3.551402e+03)*S24+(-1.033039e+01)*S25+(-2.834998e+00)*S26+2.603831e+02*S27+(-4.974715e+00)*S28+(-2.510424e+01)*S29'
.param V3_part4='V3_part3+(-5.875107e+01)*S30+(-2.948945e+01)*S31+(-9.774699e+00)*S32+1.441091e+02*S33+(-3.939830e+00)*S34+(-4.498863e+00)*S35+(-8.603012e+00)*S36+(-7.053222e+00)*S37+(-1.499379e+01)*S38+(-3.004890e-02)*S39'
.param V3='V3_part4+(-2.491473e+00)*S40+(-2.264026e+01)*S41+(-5.140598e-01)*S42+(-7.670072e+00)*S43+(-1.333403e+01)*S44'
.param V4_part1='2.419937e+00*S0+1.241373e+00*S1+1.018107e+03*S2+4.514560e+02*S3+1.942794e+00*S4+1.182359e+00*S5+1.801469e+00*S6+1.369358e+03*S7+1.451777e+00*S8+2.425858e+02*S9'
.param V4_part2='V4_part1+1.447778e+00*S10+8.816683e-01*S11+3.621733e+00*S12+3.140416e+00*S13+3.025460e+00*S14+1.045934e+03*S15+1.399677e+00*S16+(-3.593073e+02)*S17+2.748045e+02*S18+2.246901e+00*S19'
.param V4_part3='V4_part2+1.339032e+00*S20+3.963271e+00*S21+4.731523e+03*S22+3.464887e+00*S23+1.000000e+04*S24+8.134977e+02*S25+2.389341e+00*S26+3.660988e+03*S27+3.325062e+01*S28+5.761678e+01*S29'
.param V4_part4='V4_part3+2.293023e+03*S30+1.694367e+02*S31+2.180847e+01*S32+5.127028e+03*S33+1.682515e+01*S34+4.782988e+00*S35+5.715569e+01*S36+2.844161e+01*S37+3.587996e+01*S38+2.716898e+01*S39'
.param V4='V4_part4+5.969831e+00*S40+4.497173e+01*S41+4.689245e-01*S42+3.821804e+01*S43+3.439074e+01*S44'
.param V5_part1='3.654794e-01*S0+4.367595e-01*S1+(-3.805465e+01)*S2+4.708471e+02*S3+9.669987e-01*S4+8.969552e-01*S5+2.435514e-01*S6+5.153985e+02*S7+4.562221e-01*S8+1.141878e+02*S9'
.param V5_part2='V5_part1+6.769870e-01*S10+6.532968e-01*S11+5.206846e-01*S12+9.683459e-01*S13+1.372975e+00*S14+3.618500e+02*S15+4.693173e-01*S16+5.485121e+02*S17+2.491786e+02*S18+1.094949e+00*S19'
.param V5_part3='V5_part2+1.016113e+00*S20+7.523114e-01*S21+(-4.429492e+02)*S22+3.398039e+00*S23+1.106716e+03*S24+(-5.634158e+01)*S25+2.975483e+00*S26+(-1.467912e+02)*S27+1.114588e+00*S28+3.411129e+00*S29'
.param V5_part4='V5_part3+(-4.606212e+01)*S30+(-1.936245e+00)*S31+2.115924e+00*S32+(-1.609182e+02)*S33+1.649797e+00*S34+4.711860e+00*S35+1.603745e+00*S36+1.648784e+00*S37+2.959845e+00*S38+9.937261e-01*S39'
.param V5='V5_part4+2.542665e+00*S40+3.604157e+00*S41+4.092008e+00*S42+2.060539e+00*S43+3.647729e+00*S44'
.param V6_part1='(-1.521770e-02)*S0+(-1.790041e-02)*S1+0.000000e+00*S2+(-1.065910e+00)*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+3.695703e+00*S7+(-3.767940e-02)*S8+0.000000e+00*S9'
.param V6_part2='V6_part1+0.000000e+00*S10+(-2.816604e-02)*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+1.601405e+00*S15+2.940280e-02*S16+0.000000e+00*S17+(-7.258362e-01)*S18+0.000000e+00*S19'
.param V6_part3='V6_part2+0.000000e+00*S20+0.000000e+00*S21+(-8.253207e+00)*S22+0.000000e+00*S23+9.525422e-02*S24+0.000000e+00*S25+0.000000e+00*S26+(-2.673879e+00)*S27+1.537487e-01*S28+1.844659e-01*S29'
.param V6_part4='V6_part3+0.000000e+00*S30+0.000000e+00*S31+(-1.357696e+00)*S32+(-3.325824e+00)*S33+(-8.331566e-03)*S34+0.000000e+00*S35+4.409937e-02*S36+(-2.170019e-01)*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V6='V6_part4+2.047468e-01*S40+0.000000e+00*S41+(-1.221960e-02)*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V7_part1='1.160475e-01*S0+5.813486e-02*S1+0.000000e+00*S2+5.749401e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+7.039274e+00*S7+5.477436e-02*S8+0.000000e+00*S9'
.param V7_part2='V7_part1+0.000000e+00*S10+4.790836e-02*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+8.623488e+00*S15+1.815293e-01*S16+0.000000e+00*S17+2.066741e+00*S18+0.000000e+00*S19'
.param V7_part3='V7_part2+0.000000e+00*S20+0.000000e+00*S21+1.894503e+01*S22+0.000000e+00*S23+5.379948e+01*S24+0.000000e+00*S25+0.000000e+00*S26+1.761732e+01*S27+(-2.792273e-01)*S28+1.594073e-01*S29'
.param V7_part4='V7_part3+0.000000e+00*S30+0.000000e+00*S31+2.698570e+00*S32+4.787549e+01*S33+2.445747e-01*S34+0.000000e+00*S35+2.375024e-02*S36+3.878740e-01*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V7='V7_part4+(-1.746093e-01)*S40+0.000000e+00*S41+1.783805e-01*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V8_part1='2.522983e-02*S0+(-2.242802e-03)*S1+0.000000e+00*S2+4.146170e-01*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+(-3.737858e+00)*S7+6.953769e-03*S8+0.000000e+00*S9'
.param V8_part2='V8_part1+0.000000e+00*S10+1.541927e-02*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+(-3.439341e+00)*S15+2.730651e-02*S16+0.000000e+00*S17+6.420549e-01*S18+0.000000e+00*S19'
.param V8_part3='V8_part2+0.000000e+00*S20+0.000000e+00*S21+9.360077e+00*S22+0.000000e+00*S23+(-1.654555e+01)*S24+0.000000e+00*S25+0.000000e+00*S26+2.515257e+00*S27+4.241821e-01*S28+(-1.059681e-01)*S29'
.param V8_part4='V8_part3+0.000000e+00*S30+0.000000e+00*S31+(-5.474835e-01)*S32+(-4.220350e+00)*S33+4.089720e-01*S34+0.000000e+00*S35+1.559584e-01*S36+7.838251e-01*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V8='V8_part4+1.743153e-02*S40+0.000000e+00*S41+1.847904e-01*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V9_part1='(-9.972657e-02)*S0+8.142120e-02*S1+0.000000e+00*S2+1.443367e+02*S3+(-6.927764e-02)*S4+9.393997e-02*S5+(-2.241444e-01)*S6+0.000000e+00*S7+(-1.802346e-01)*S8+0.000000e+00*S9'
.param V9_part2='V9_part1+(-1.834675e-01)*S10+(-3.594864e-02)*S11+(-1.479409e-01)*S12+(-1.864345e-01)*S13+(-2.290860e-01)*S14+0.000000e+00*S15+6.130910e-02*S16+0.000000e+00*S17+0.000000e+00*S18+(-1.034067e-01)*S19'
.param V9_part3='V9_part2+9.972946e-02*S20+2.622105e-02*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+(-2.684448e+00)*S28+0.000000e+00*S29'
.param V9_part4='V9_part3+0.000000e+00*S30+0.000000e+00*S31+(-1.191368e+01)*S32+0.000000e+00*S33+(-1.330708e+00)*S34+0.000000e+00*S35+2.425748e+00*S36+(-4.914357e+00)*S37+(-1.999638e+01)*S38+6.339533e-02*S39'
.param V9='V9_part4+(-1.085301e-01)*S40+(-1.216801e+01)*S41+0.000000e+00*S42+(-5.407233e+00)*S43+(-1.667380e+01)*S44'
.param V10_part1='(-3.650109e-02)*S0+8.258838e-02*S1+0.000000e+00*S2+(-2.125153e+01)*S3+1.583079e-03*S4+1.695513e-02*S5+(-7.288176e-02)*S6+0.000000e+00*S7+(-5.295038e-02)*S8+0.000000e+00*S9'
.param V10_part2='V10_part1+(-4.959436e-02)*S10+2.048416e-02*S11+3.931349e-02*S12+9.560010e-02*S13+5.852672e-02*S14+0.000000e+00*S15+1.510254e-01*S16+0.000000e+00*S17+0.000000e+00*S18+5.589892e-03*S19'
.param V10_part3='V10_part2+2.887384e-02*S20+(-1.111410e-01)*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+7.198464e+01*S28+0.000000e+00*S29'
.param V10_part4='V10_part3+0.000000e+00*S30+0.000000e+00*S31+2.247178e+01*S32+0.000000e+00*S33+6.413825e+00*S34+0.000000e+00*S35+(-6.933581e+00)*S36+2.479737e+01*S37+5.525695e+01*S38+1.974621e+01*S39'
.param V10='V10_part4+1.611263e-01*S40+2.655706e+01*S41+0.000000e+00*S42+7.682372e+01*S43+5.906140e+01*S44'
.param V11_part1='2.864114e-01*S0+1.866587e-01*S1+0.000000e+00*S2+(-6.869345e+01)*S3+2.882013e-01*S4+1.849317e-01*S5+2.568509e-01*S6+0.000000e+00*S7+2.382855e-01*S8+0.000000e+00*S9'
.param V11_part2='V11_part1+2.443039e-01*S10+1.358670e-01*S11+3.000288e-01*S12+2.917959e-01*S13+3.315428e-01*S14+0.000000e+00*S15+1.895269e-01*S16+0.000000e+00*S17+0.000000e+00*S18+2.978714e-01*S19'
.param V11_part3='V11_part2+1.879347e-01*S20+3.748971e-01*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+(-2.766016e+00)*S28+0.000000e+00*S29'
.param V11_part4='V11_part3+0.000000e+00*S30+0.000000e+00*S31+7.530563e-01*S32+0.000000e+00*S33+5.799913e-01*S34+0.000000e+00*S35+2.946493e-01*S36+4.973405e-01*S37+(-1.002327e+00)*S38+4.196765e-01*S39'
.param V11='V11_part4+4.926273e-01*S40+7.326007e-01*S41+0.000000e+00*S42+(-2.563881e+00)*S43+(-1.732824e+00)*S44'
.param V12_part1='(-4.107151e-01)*S0+1.009052e+00*S1+5.598906e-02*S2+2.460860e-02*S3+(-3.945829e+01)*S4+7.012444e+00*S5+1.921148e+00*S6+(-3.281457e-03)*S7+(-1.307818e+02)*S8+(-2.548270e-03)*S9'
.param V12_part2='V12_part1+(-4.512403e+02)*S10+1.208097e+01*S11+1.592168e+00*S12+(-3.985514e+01)*S13+(-1.573979e+02)*S14+(-1.360479e-02)*S15+3.387694e-01*S16+(-5.212354e-03)*S17+5.281665e-02*S18+(-5.907660e+01)*S19'
.param V12_part3='V12_part2+6.553917e+00*S20+(-1.428040e+00)*S21+8.247486e-02*S22+(-5.579239e+00)*S23+(-1.708872e-02)*S24+9.236705e-02*S25+(-3.689253e+00)*S26+5.593763e-02*S27+7.302127e-01*S28+1.128619e+00*S29'
.param V12_part4='V12_part3+5.356814e-02*S30+3.042044e-01*S31+2.001160e+00*S32+5.773848e-02*S33+3.460359e+00*S34+(-1.122587e+01)*S35+2.104932e-01*S36+1.001945e+00*S37+1.954837e+00*S38+1.185788e+00*S39'
.param V12='V12_part4+(-5.146991e+01)*S40+3.870168e+00*S41+(-6.830589e-01)*S42+1.183579e+00*S43+3.997558e+00*S44'
.param V13_part1='4.971914e+01*S0+1.844183e+01*S1+1.078316e+00*S2+9.533224e-01*S3+7.971047e+01*S4+7.144990e+01*S5+3.692285e+01*S6+5.513354e-01*S7+9.064488e+02*S8+6.318470e-01*S9'
.param V13_part2='V13_part1+1.179988e+03*S10+1.139216e+02*S11+7.116204e+01*S12+1.681909e+02*S13+2.658751e+02*S14+1.158615e+00*S15+1.385418e+01*S16+1.433044e+00*S17+1.167455e+00*S18+1.241126e+02*S19'
.param V13_part3='V13_part2+5.302835e+01*S20+2.500439e+01*S21+2.814720e+00*S22+1.499576e+01*S23+2.003467e+00*S24+2.235300e+00*S25+9.719817e+00*S26+3.666364e+00*S27+4.820750e+00*S28+4.495241e+00*S29'
.param V13_part4='V13_part3+3.020985e+00*S30+3.632932e+00*S31+3.971694e+00*S32+4.680070e+00*S33+9.234622e+00*S34+2.962977e+01*S35+5.911682e+00*S36+5.982325e+00*S37+4.954659e+00*S38+9.190408e+00*S39'
.param V13='V13_part4+1.406444e+02*S40+8.217888e+00*S41+1.073310e+01*S42+7.268852e+00*S43+5.472518e+00*S44'
.param V14_part1='(-9.025067e+00)*S0+(-3.373727e+00)*S1+(-1.604021e-01)*S2+(-2.738216e-02)*S3+1.760145e+00*S4+(-3.426070e+01)*S5+(-1.000808e+01)*S6+(-3.652044e-03)*S7+1.527110e+02*S8+(-4.049058e-02)*S9'
.param V14_part2='V14_part1+4.970059e+02*S10+(-2.701087e+01)*S11+(-2.037368e+01)*S12+8.378409e+00*S13+1.099365e+02*S14+(-2.780821e-02)*S15+(-2.090528e+00)*S16+(-9.734171e-02)*S17+(-5.549156e-02)*S18+(-3.484951e-02)*S19'
.param V14_part3='V14_part2+(-2.636141e+01)*S20+(-1.724910e+00)*S21+(-2.608135e-01)*S22+2.622665e-01*S23+5.696241e-02*S24+(-3.012770e-01)*S25+2.160149e+00*S26+1.866324e-01*S27+(-9.674446e-01)*S28+(-1.831747e+00)*S29'
.param V14_part4='V14_part3+9.657547e-02*S30+(-8.160525e-01)*S31+(-2.026105e+00)*S32+3.913144e-01*S33+(-5.494656e+00)*S34+3.578345e+00*S35+(-4.055522e-01)*S36+(-2.003313e+00)*S37+(-1.883170e+00)*S38+7.895323e-01*S39'
.param V14='V14_part4+7.496281e+01*S40+(-5.596417e+00)*S41+2.408947e+00*S42+(-1.287358e+00)*S43+(-2.347544e+00)*S44'
.param V15_part1='(-3.330399e+02)*S0+(-1.056029e+02)*S1+(-8.472364e-01)*S2+(-4.412290e-01)*S3+(-5.757349e+02)*S4+(-1.130645e+03)*S5+(-4.263397e+02)*S6+(-1.914478e-01)*S7+1.000000e+04*S8+(-3.394309e-01)*S9'
.param V15_part2='V15_part1+1.000000e+04*S10+1.357549e+02*S11+(-5.868757e+02)*S12+(-2.508688e+02)*S13+(-1.595201e+03)*S14+(-4.355533e-01)*S15+(-4.091731e+01)*S16+(-8.799458e-01)*S17+(-4.269780e-01)*S18+(-8.972050e+02)*S19'
.param V15_part3='V15_part2+(-5.152304e+02)*S20+(-3.515772e+01)*S21+(-1.614133e+00)*S22+(-9.923818e+00)*S23+(-5.830611e-01)*S24+(-1.600829e+00)*S25+(-1.208075e+01)*S26+(-6.366037e-01)*S27+(-2.815315e+00)*S28+(-4.034188e+00)*S29'
.param V15_part4='V15_part3+(-6.243476e-01)*S30+(-1.256277e+00)*S31+(-3.843396e+00)*S32+(-6.076530e-01)*S33+(-4.168426e+00)*S34+(-1.391710e+01)*S35+7.187790e-01*S36+(-2.958361e+00)*S37+(-4.562121e+00)*S38+(-1.629376e+00)*S39'
.param V15='V15_part4+(-2.596253e+01)*S40+(-3.029031e+00)*S41+(-2.072831e+00)*S42+(-2.956431e+00)*S43+(-5.668712e+00)*S44'
.param V16_part1='8.139260e+02*S0+1.954515e+02*S1+1.866585e+00*S2+1.181649e+00*S3+1.463636e+03*S4+9.299449e+02*S5+9.352280e+02*S6+9.983200e-01*S7+8.381181e+03*S8+8.456443e-01*S9'
.param V16_part2='V16_part1+8.968823e+03*S10+1.144681e+03*S11+1.390069e+03*S12+6.116138e+03*S13+5.518699e+03*S14+2.768135e+00*S15+1.121167e+02*S16+2.209189e+00*S17+1.326889e+00*S18+2.362535e+03*S19'
.param V16_part3='V16_part2+3.579237e+02*S20+5.998067e+02*S21+3.885939e+00*S22+2.395790e+01*S23+4.166761e+00*S24+3.256695e+00*S25+2.386342e+01*S26+5.080870e+00*S27+4.583540e+00*S28+4.300026e+00*S29'
.param V16_part4='V16_part3+4.471680e+00*S30+3.087226e+00*S31+2.794545e+00*S32+5.981621e+00*S33+1.714044e+00*S34+3.483109e+01*S35+1.564473e-01*S36+4.132931e+00*S37+4.697114e+00*S38+2.908129e+00*S39'
.param V16='V16_part4+4.131345e+02*S40+2.713855e+00*S41+2.593408e+01*S42+5.475887e+00*S43+6.119903e+00*S44'
.param V17_part1='3.160653e+02*S0+1.281472e+02*S1+6.693667e-01*S2+6.398810e-01*S3+(-7.042891e+01)*S4+1.018601e+03*S5+2.401482e+02*S6+2.925906e-01*S7+1.000000e+04*S8+4.512834e-01*S9'
.param V17_part2='V17_part1+1.000000e+04*S10+8.721360e+02*S11+2.791583e+02*S12+(-4.400006e+02)*S13+(-4.392228e+02)*S14+4.029960e-01*S15+8.066389e+01*S16+7.117274e-01*S17+6.873448e-01*S18+(-1.366961e+02)*S19'
.param V17_part3='V17_part2+5.647541e+02*S20+(-3.587675e+00)*S21+1.243474e+00*S22+2.045644e+00*S23+5.612280e-01*S24+1.127154e+00*S25+1.675851e+00*S26+9.352159e-01*S27+2.893501e+00*S28+3.294920e+00*S29'
.param V17_part4='V17_part3+8.052384e-01*S30+1.550082e+00*S31+4.250039e+00*S32+1.134998e+00*S33+7.423126e+00*S34+3.287898e+00*S35+1.824024e+00*S36+3.694817e+00*S37+4.072799e+00*S38+4.341567e+00*S39'
.param V17='V17_part4+(-1.736554e+01)*S40+6.163497e+00*S41+1.105165e+00*S42+3.667667e+00*S43+4.921686e+00*S44'
.param V18_part1='1.140212e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-4.630095e-02)*S3+0.000000e+00*S4+1.146342e+00*S5+1.057392e+00*S6+(-7.567239e-03)*S7+1.894912e+01*S8+0.000000e+00*S9'
.param V18_part2='V18_part1+(-1.581908e+02)*S10+(-3.557346e+00)*S11+0.000000e+00*S12+(-9.469270e+00)*S13+0.000000e+00*S14+2.550944e-02*S15+6.160488e-01*S16+0.000000e+00*S17+(-5.017651e-02)*S18+0.000000e+00*S19'
.param V18_part3='V18_part2+0.000000e+00*S20+0.000000e+00*S21+7.219413e-05*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+(-2.085876e-01)*S26+0.000000e+00*S27+0.000000e+00*S28+2.866226e-01*S29'
.param V18_part4='V18_part3+0.000000e+00*S30+0.000000e+00*S31+(-1.024472e-01)*S32+7.034574e-02*S33+0.000000e+00*S34+0.000000e+00*S35+6.031298e-02*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V18='V18_part4+0.000000e+00*S40+(-2.066786e-01)*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V19_part1='7.534808e+00*S0+0.000000e+00*S1+0.000000e+00*S2+1.033342e-01*S3+0.000000e+00*S4+1.083709e+01*S5+1.413420e+00*S6+5.960615e-02*S7+3.510867e+02*S8+0.000000e+00*S9'
.param V19_part2='V19_part1+4.306731e+02*S10+2.259065e+01*S11+0.000000e+00*S12+3.448186e+01*S13+0.000000e+00*S14+1.363307e-01*S15+8.314068e-01*S16+0.000000e+00*S17+1.666385e-01*S18+0.000000e+00*S19'
.param V19_part3='V19_part2+0.000000e+00*S20+0.000000e+00*S21+1.196260e-01*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+3.772036e-01*S26+0.000000e+00*S27+0.000000e+00*S28+(-3.087033e-02)*S29'
.param V19_part4='V19_part3+0.000000e+00*S30+0.000000e+00*S31+3.520711e-01*S32+1.216768e-01*S33+0.000000e+00*S34+0.000000e+00*S35+(-1.226415e-01)*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V19='V19_part4+0.000000e+00*S40+2.680457e-01*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V20_part1='(-2.248132e+00)*S0+0.000000e+00*S1+0.000000e+00*S2+4.866208e-03*S3+0.000000e+00*S4+(-5.482758e+00)*S5+(-1.999934e+00)*S6+(-1.465027e-02)*S7+(-7.014033e+01)*S8+0.000000e+00*S9'
.param V20_part2='V20_part1+4.160583e+01*S10+(-1.687613e+00)*S11+0.000000e+00*S12+6.983120e+00*S13+0.000000e+00*S14+2.253388e-02*S15+(-2.421554e-01)*S16+0.000000e+00*S17+4.110136e-02*S18+0.000000e+00*S19'
.param V20_part3='V20_part2+0.000000e+00*S20+0.000000e+00*S21+(-8.098463e-02)*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+3.485960e-01*S26+0.000000e+00*S27+0.000000e+00*S28+1.764632e-01*S29'
.param V20_part4='V20_part3+0.000000e+00*S30+0.000000e+00*S31+5.419639e-02*S32+(-2.364371e-02)*S33+0.000000e+00*S34+0.000000e+00*S35+(-2.022397e-04)*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V20='V20_part4+0.000000e+00*S40+4.479457e-02*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V21_part1='0.000000e+00*S0+0.000000e+00*S1+(-1.151104e-01)*S2+9.807137e-02*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+(-3.945254e-02)*S7+0.000000e+00*S8+(-3.133941e-02)*S9'
.param V21_part2='V21_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+(-1.173709e-01)*S15+0.000000e+00*S16+(-1.230967e-01)*S17+4.971823e-02*S18+0.000000e+00*S19'
.param V21_part3='V21_part2+0.000000e+00*S20+0.000000e+00*S21+(-1.247222e-01)*S22+(-1.467708e+01)*S23+(-1.490234e-01)*S24+(-2.302528e-01)*S25+(-1.302288e+01)*S26+(-3.882734e-02)*S27+0.000000e+00*S28+(-1.572562e-01)*S29'
.param V21_part4='V21_part3+(-4.770668e-02)*S30+(-5.363986e-01)*S31+0.000000e+00*S32+1.107176e-01*S33+0.000000e+00*S34+(-2.272573e+01)*S35+(-9.128305e-01)*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V21='V21_part4+0.000000e+00*S40+0.000000e+00*S41+(-2.463903e-01)*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V22_part1='0.000000e+00*S0+0.000000e+00*S1+8.486070e-02*S2+3.885823e-02*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+8.931019e-03*S7+0.000000e+00*S8+3.222737e-02*S9'
.param V22_part2='V22_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+1.551432e-02*S15+0.000000e+00*S16+5.691755e-02*S17+8.016420e-02*S18+0.000000e+00*S19'
.param V22_part3='V22_part2+0.000000e+00*S20+0.000000e+00*S21+1.024767e-01*S22+3.817748e+01*S23+(-3.278056e-02)*S24+1.228049e-01*S25+2.178192e+01*S26+2.265291e-02*S27+0.000000e+00*S28+(-4.784756e-01)*S29'
.param V22_part4='V22_part3+(-1.116167e-02)*S30+2.418515e-01*S31+0.000000e+00*S32+1.215247e-01*S33+0.000000e+00*S34+5.810043e+01*S35+7.829885e-01*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V22='V22_part4+0.000000e+00*S40+0.000000e+00*S41+1.507747e+01*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V23_part1='0.000000e+00*S0+0.000000e+00*S1+2.848087e-01*S2+1.789799e-01*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+1.445741e-01*S7+0.000000e+00*S8+1.361638e-01*S9'
.param V23_part2='V23_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+2.873356e-01*S15+0.000000e+00*S16+2.839914e-01*S17+2.037815e-01*S18+0.000000e+00*S19'
.param V23_part3='V23_part2+0.000000e+00*S20+0.000000e+00*S21+3.731026e-01*S22+(-2.183328e-02)*S23+2.977657e-01*S24+3.250646e-01*S25+1.416822e+00*S26+3.588132e-01*S27+0.000000e+00*S28+8.001163e-01*S29'
.param V23_part4='V23_part3+3.681209e-01*S30+5.639708e-01*S31+0.000000e+00*S32+3.801027e-01*S33+0.000000e+00*S34+(-7.008157e-01)*S35+8.565091e-01*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V23='V23_part4+0.000000e+00*S40+0.000000e+00*S41+5.336401e-01*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V24_part1='1.238894e+00*S0+1.228651e+00*S1+1.716420e+00*S2+1.135736e+00*S3+2.046361e+00*S4+1.386666e+00*S5+1.504166e+00*S6+9.851368e-01*S7+1.135250e+00*S8+1.509744e+00*S9'
.param V24_part2='V24_part1+1.497971e+00*S10+1.230426e+00*S11+1.601729e+00*S12+1.779394e+00*S13+2.585868e+00*S14+2.501201e+00*S15+8.334163e+00*S16+1.543282e+00*S17+9.744565e-01*S18+2.022939e+00*S19'
.param V24_part3='V24_part2+1.446739e+00*S20+(-7.074039e+00)*S21+2.823049e+00*S22+5.939577e+00*S23+1.622803e+00*S24+3.039278e+00*S25+5.736007e+01*S26+2.409325e+00*S27+4.619249e+00*S28+1.144747e+02*S29'
.param V24_part4='V24_part3+2.277301e+00*S30+4.299893e-01*S31+3.764883e+00*S32+4.052168e+00*S33+1.029031e+02*S34+5.184533e+00*S35+6.250000e+02*S36+4.336765e+02*S37+5.540744e+00*S38+3.722151e+00*S39'
.param V24='V24_part4+8.459561e+00*S40+7.972298e+03*S41+1.622698e+01*S42+5.712886e+00*S43+9.476562e+00*S44'
.param V25_part1='2.211609e+00*S0+1.231666e+00*S1+4.095931e-01*S2+9.832169e-01*S3+1.336013e-01*S4+2.594167e-01*S5+3.136187e-01*S6+1.196734e+00*S7+3.729888e-01*S8+2.184456e-01*S9'
.param V25_part2='V25_part1+3.622352e-02*S10+3.632140e-01*S11+1.468828e+00*S12+8.934856e-01*S13+3.621739e-01*S14+1.277970e+00*S15+(-2.254776e+00)*S16+7.305313e-01*S17+1.771752e+00*S18+7.562926e-02*S19'
.param V25_part3='V25_part2+3.562430e-01*S20+2.279408e+01*S21+1.712775e+00*S22+2.056084e+00*S23+1.307896e+00*S24+1.724720e+00*S25+4.438233e+03*S26+1.916153e+00*S27+4.379878e+00*S28+(-6.533702e+01)*S29'
.param V25_part4='V25_part3+1.363187e+00*S30+8.500078e+00*S31+4.754973e+00*S32+2.630560e+00*S33+2.147337e+03*S34+3.961687e+00*S35+1.000000e+04*S36+3.777675e+03*S37+3.724268e+00*S38+8.113474e+00*S39'
.param V25='V25_part4+2.129203e+00*S40+5.549391e+03*S41+2.025796e+01*S42+3.444703e+00*S43+1.242782e+00*S44'
.param V26_part1='(-5.436294e-01)*S0+(-2.782261e-01)*S1+(-5.432445e-01)*S2+(-3.543316e-01)*S3+(-7.362981e-01)*S4+(-2.611828e-01)*S5+(-4.536893e-01)*S6+(-3.598207e-01)*S7+(-5.151540e-01)*S8+(-2.871186e-01)*S9'
.param V26_part2='V26_part1+(-6.375622e-01)*S10+(-2.139400e-01)*S11+(-7.623068e-01)*S12+(-1.293135e+00)*S13+(-1.679389e+00)*S14+(-7.985440e-01)*S15+1.188477e+00*S16+(-8.618175e-01)*S17+8.201219e-02*S18+(-7.701689e-01)*S19'
.param V26_part3='V26_part2+(-2.323714e-01)*S20+7.594332e+01*S21+(-3.028334e+00)*S22+(-6.369508e+00)*S23+(-9.129083e-01)*S24+(-2.973508e+00)*S25+(-1.280322e+00)*S26+(-1.906727e+00)*S27+(-6.271298e+00)*S28+(-2.589260e+01)*S29'
.param V26_part4='V26_part3+(-1.479683e+00)*S30+4.492150e+00*S31+(-3.419323e+00)*S32+(-3.833237e+00)*S33+1.657996e+02*S34+(-6.326594e+00)*S35+1.000000e+04*S36+3.869737e+03*S37+(-7.328498e+00)*S38+(-2.221043e+00)*S39'
.param V26='V26_part4+(-1.017392e+01)*S40+4.475144e+03*S41+4.573612e+00*S42+(-6.203764e+00)*S43+(-9.624129e+00)*S44'
.param V27_part1='(-1.062322e+00)*S0+1.648113e+00*S1+1.958236e+00*S2+6.958703e-01*S3+1.846024e+00*S4+3.331497e+00*S5+5.368994e+00*S6+8.879146e+00*S7+(-8.652594e+00)*S8+3.180758e+00*S9'
.param V27_part2='V27_part1+1.836793e+00*S10+(-2.722433e+00)*S11+2.374310e+00*S12+2.663435e+00*S13+1.412887e+00*S14+3.217994e+01*S15+2.522098e+01*S16+1.930317e+00*S17+3.548817e-01*S18+1.567720e+00*S19'
.param V27_part3='V27_part2+2.146023e+00*S20+1.944436e+00*S21+5.494765e-03*S22+3.202691e+00*S23+8.832351e+00*S24+2.842151e+00*S25+3.926568e+00*S26+1.668100e+00*S27+3.293964e+00*S28+1.320559e+01*S29'
.param V27_part4='V27_part3+1.523827e+00*S30+3.035126e+00*S31+(-3.428735e+00)*S32+(-1.562367e+02)*S33+6.935532e+00*S34+4.721654e+00*S35+4.754522e+00*S36+4.681608e+00*S37+4.574558e+00*S38+2.747858e+00*S39'
.param V27='V27_part4+8.787670e+00*S40+4.709881e+00*S41+1.675871e+00*S42+2.911410e+00*S43+4.798850e+00*S44'
.param V28_part1='1.667495e+01*S0+2.657517e+00*S1+1.152758e+00*S2+5.044444e+00*S3+9.914982e-01*S4+1.273979e+00*S5+(-2.194869e+00)*S6+1.782940e+00*S7+2.705315e+01*S8+3.853638e-01*S9'
.param V28_part2='V28_part1+5.163303e+00*S10+8.348056e+00*S11+3.818652e+00*S12+1.920988e+00*S13+2.292481e+00*S14+(-2.308180e+01)*S15+(-1.957817e-01)*S16+7.735034e-01*S17+4.843828e+00*S18+9.288786e-01*S19'
.param V28_part3='V28_part2+7.716093e-01*S20+1.226299e+00*S21+1.130114e+01*S22+5.168390e-01*S23+8.553918e+00*S24+9.404816e-01*S25+1.227963e-01*S26+7.365877e+00*S27+1.092175e+00*S28+(-6.113150e+00)*S29'
.param V28_part4='V28_part3+4.666634e+00*S30+5.744979e-01*S31+1.409890e+01*S32+2.467260e+03*S33+2.928080e-01*S34+7.002255e-01*S35+5.019258e-04*S36+9.486107e-01*S37+5.773953e-01*S38+4.727704e+00*S39'
.param V28='V28_part4+(-4.592397e+00)*S40+1.730745e+00*S41+6.286523e+00*S42+2.603017e+00*S43+4.323968e-02*S44'
.param V29_part1='6.907880e+00*S0+(-4.737251e-01)*S1+1.739703e-01*S2+4.207026e-01*S3+5.224602e-01*S4+(-6.201496e-01)*S5+(-1.414645e+00)*S6+(-4.883219e+00)*S7+1.948278e+01*S8+(-2.198082e-01)*S9'
.param V29_part2='V29_part1+6.255391e+00*S10+6.343953e+00*S11+(-1.399942e+00)*S12+3.608723e+00*S13+2.114948e+00*S14+(-1.542124e+01)*S15+(-1.633732e+01)*S16+(-8.040823e-02)*S17+4.716302e-01*S18+2.912389e-01*S19'
.param V29_part3='V29_part2+(-4.956964e-01)*S20+(-1.519238e+00)*S21+1.652734e+00*S22+3.282940e-01*S23+(-5.012517e+00)*S24+1.751417e+00*S25+(-2.667420e+00)*S26+2.531945e+00*S27+5.669585e-01*S28+4.807435e+00*S29'
.param V29_part4='V29_part3+2.376308e-01*S30+(-2.335347e+00)*S31+(-3.336156e+00)*S32+1.219551e+03*S33+(-4.903618e+00)*S34+(-6.278267e-01)*S35+(-2.822982e+00)*S36+(-3.671629e+00)*S37+2.220184e-01*S38+(-4.917330e-01)*S39'
.param V29='V29_part4+1.874539e+00*S40+(-3.674897e+00)*S41+1.262490e-01*S42+(-2.533921e-01)*S43+(-1.171375e-02)*S44'
.param V30_part1='(-2.008183e+00)*S0+1.134886e+01*S1+(-3.271509e+01)*S2+1.662765e+00*S3+(-4.515517e+01)*S4+1.104234e+01*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V30_part2='V30_part1+1.774053e+01*S10+0.000000e+00*S11+(-1.815412e+00)*S12+(-2.805312e+01)*S13+(-1.538184e+01)*S14+1.254477e+00*S15+(-4.293105e+00)*S16+5.050786e+00*S17+(-3.235690e+00)*S18+(-5.179061e+01)*S19'
.param V30_part3='V30_part2+8.381790e+00*S20+(-4.667734e+00)*S21+(-1.089658e+01)*S22+7.229578e+01*S23+(-4.042523e+00)*S24+0.000000e+00*S25+(-7.242943e+00)*S26+(-2.983054e+01)*S27+4.535324e+00*S28+2.457131e+01*S29'
.param V30_part4='V30_part3+(-2.652386e+01)*S30+(-2.228350e+01)*S31+(-2.280133e+01)*S32+(-8.570364e+00)*S33+(-2.954098e+01)*S34+3.686670e+01*S35+(-2.481519e+00)*S36+(-1.389928e+01)*S37+4.683298e+01*S38+8.749116e+00*S39'
.param V30='V30_part4+(-7.261285e+01)*S40+6.545808e+01*S41+1.446734e+01*S42+(-2.242695e+01)*S43+(-6.576940e+01)*S44'
.param V31_part1='2.931256e+01*S0+3.134386e+01*S1+6.578100e+01*S2+3.606056e+01*S3+6.731886e+01*S4+3.313756e+01*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V31_part2='V31_part1+(-5.748989e+00)*S10+0.000000e+00*S11+7.849761e+01*S12+8.601448e+01*S13+8.611795e+01*S14+3.458332e+01*S15+6.902161e+01*S16+1.809711e+01*S17+7.904986e+01*S18+9.171555e+01*S19'
.param V31_part3='V31_part2+3.998371e+01*S20+1.183244e+02*S21+1.187315e+02*S22+(-1.787946e+01)*S23+9.991959e+01*S24+0.000000e+00*S25+8.576182e+01*S26+1.531126e+02*S27+9.304424e+01*S28+1.296847e+01*S29'
.param V31_part4='V31_part3+1.505163e+02*S30+1.567081e+02*S31+1.454677e+02*S32+1.866792e+02*S33+1.967937e+02*S34+1.143362e+02*S35+1.035788e+02*S36+1.619033e+02*S37+2.529944e+01*S38+2.020457e+02*S39'
.param V31='V31_part4+1.236838e+02*S40+1.437279e+02*S41+1.697528e+02*S42+2.040266e+02*S43+2.317936e+02*S44'
.param V32_part1='7.432665e+00*S0+(-9.573129e+00)*S1+3.198080e+01*S2+2.537770e+00*S3+3.283990e+01*S4+(-6.590024e+00)*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V32_part2='V32_part1+(-1.352770e+01)*S10+0.000000e+00*S11+2.916038e+01*S12+3.465804e+01*S13+3.952301e+01*S14+1.111942e+01*S15+6.384424e+00*S16+2.537699e+01*S17+(-5.226532e+00)*S18+2.844104e+01*S19'
.param V32_part3='V32_part2+1.560793e+01*S20+4.076935e+01*S21+4.907144e+01*S22+4.030711e+01*S23+2.496857e+01*S24+0.000000e+00*S25+3.533191e+01*S26+9.843828e+01*S27+1.664446e+01*S28+1.506708e+02*S29'
.param V32_part4='V32_part3+7.041601e+01*S30+(-2.289991e+01)*S31+(-8.229941e+01)*S32+8.209232e+01*S33+1.173482e+02*S34+7.147002e+00*S35+5.933112e+01*S36+7.229457e+01*S37+1.276807e+02*S38+3.319652e+01*S39'
.param V32='V32_part4+3.119837e+02*S40+(-1.260382e+02)*S41+2.536682e+00*S42+1.084209e+02*S43+1.445793e+02*S44'
.param V33_part1='0.000000e+00*S0+(-1.773851e+01)*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+(-3.293577e+01)*S5+0.000000e+00*S6+(-1.497692e+01)*S7+0.000000e+00*S8+(-1.684053e+01)*S9'
.param V33_part2='V33_part1+(-2.087840e+01)*S10+(-4.260842e+01)*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+(-1.235929e+01)*S15+0.000000e+00*S16+(-2.528499e+01)*S17+(-8.492285e+00)*S18+0.000000e+00*S19'
.param V33_part3='V33_part2+(-4.322639e+01)*S20+0.000000e+00*S21+0.000000e+00*S22+(-1.817517e+02)*S23+0.000000e+00*S24+(-2.283381e+01)*S25+0.000000e+00*S26+4.597809e+01*S27+(-3.532472e+01)*S28+(-1.233415e+02)*S29'
.param V33_part4='V33_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+2.003890e+00*S36+0.000000e+00*S37+(-1.505676e+02)*S38+0.000000e+00*S39'
.param V33='V33_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V34_part1='0.000000e+00*S0+(-1.086712e+01)*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+1.386093e+00*S5+0.000000e+00*S6+8.250856e+01*S7+0.000000e+00*S8+6.721793e+01*S9'
.param V34_part2='V34_part1+4.534796e+01*S10+6.071422e+01*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+6.083332e+01*S15+0.000000e+00*S16+9.276250e+01*S17+(-2.740234e+01)*S18+0.000000e+00*S19'
.param V34_part3='V34_part2+4.935805e+01*S20+0.000000e+00*S21+0.000000e+00*S22+2.689817e+02*S23+0.000000e+00*S24+1.992657e+02*S25+0.000000e+00*S26+5.638995e-01*S27+1.183645e+02*S28+2.958878e+02*S29'
.param V34_part4='V34_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+9.740905e+01*S36+0.000000e+00*S37+2.769157e+02*S38+0.000000e+00*S39'
.param V34='V34_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V35_part1='0.000000e+00*S0+4.364988e+01*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+7.301274e+01*S5+0.000000e+00*S6+1.840262e+01*S7+0.000000e+00*S8+(-2.857864e+00)*S9'
.param V35_part2='V35_part1+(-1.315917e+01)*S10+1.943045e+01*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+2.029431e+01*S15+0.000000e+00*S16+(-1.044972e+01)*S17+5.735396e+01*S18+0.000000e+00*S19'
.param V35_part3='V35_part2+2.805541e+01*S20+0.000000e+00*S21+0.000000e+00*S22+2.860311e+01*S23+0.000000e+00*S24+6.302948e+01*S25+0.000000e+00*S26+(-6.707160e+01)*S27+8.827042e+01*S28+(-1.069927e+02)*S29'
.param V35_part4='V35_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-1.613676e+01)*S36+0.000000e+00*S37+(-6.326882e+01)*S38+0.000000e+00*S39'
.param V35='V35_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V36_part1='(-9.381915e-01)*S0+(-5.506246e+00)*S1+1.420258e+01*S2+(-2.996701e+00)*S3+9.229860e+00*S4+(-2.117220e+00)*S5+(-1.141332e+01)*S6+1.000000e+04*S7+(-1.065330e+00)*S8+(-1.008019e+00)*S9'
.param V36_part2='V36_part1+(-2.804059e+00)*S10+3.750979e+00*S11+(-1.724073e+02)*S12+3.731473e+00*S13+(-9.539391e+01)*S14+(-2.995600e-01)*S15+(-8.120135e-01)*S16+(-1.734455e+01)*S17+4.897796e+01*S18+1.191369e+01*S19'
.param V36_part3='V36_part2+(-1.415471e+00)*S20+(-9.464925e+00)*S21+(-5.013044e+02)*S22+(-2.000080e+03)*S23+(-2.221330e-01)*S24+(-1.999721e+03)*S25+(-2.000600e+03)*S26+(-1.998032e+03)*S27+(-1.999683e+03)*S28+(-1.332215e+02)*S29'
.param V36_part4='V36_part3+1.632393e+01*S30+1.871885e+00*S31+(-4.163311e+00)*S32+8.085403e-01*S33+2.816191e+02*S34+(-2.488680e+01)*S35+(-1.998720e+03)*S36+(-1.673783e+03)*S37+(-2.000854e+03)*S38+(-1.364405e+01)*S39'
.param V36='V36_part4+2.228570e+00*S40+(-2.281220e+01)*S41+(-2.144288e+01)*S42+(-2.417539e+02)*S43+1.799161e+02*S44'
.param V37_part1='7.942378e+00*S0+1.386566e+01*S1+1.190755e-02*S2+5.664092e+00*S3+(-9.336129e-01)*S4+5.091558e+00*S5+5.015707e+01*S6+1.000000e+04*S7+6.872481e+00*S8+2.806479e+00*S9'
.param V37_part2='V37_part1+3.043472e+00*S10+4.970212e-01*S11+9.858959e-01*S12+1.813144e-01*S13+1.190744e+00*S14+1.002361e+00*S15+(-6.402524e-01)*S16+1.197095e+00*S17+2.126497e+00*S18+(-7.648647e+00)*S19'
.param V37_part3='V37_part2+1.846331e+00*S20+(-3.852963e+00)*S21+3.603329e-01*S22+1.038777e+00*S23+4.106337e-01*S24+1.739095e+00*S25+1.730345e+00*S26+3.895647e-02*S27+9.002611e-01*S28+2.479907e+00*S29'
.param V37_part4='V37_part3+(-1.557829e+01)*S30+(-1.575340e+01)*S31+(-2.357504e+00)*S32+(-9.814811e-01)*S33+4.139231e+00*S34+2.615871e+01*S35+(-5.933580e-01)*S36+1.060160e+00*S37+2.176691e+00*S38+8.804649e+00*S39'
.param V37='V37_part4+2.306831e+01*S40+1.928455e+01*S41+1.002327e+01*S42+2.092048e+00*S43+(-1.542567e+00)*S44'
.param V38_part1='2.358973e+00*S0+6.922757e+00*S1+(-1.158863e+01)*S2+5.923717e+00*S3+(-3.799675e+00)*S4+8.405837e-01*S5+2.326803e+01*S6+1.000000e+04*S7+1.724973e+00*S8+6.379490e+00*S9'
.param V38_part2='V38_part1+7.083709e+00*S10+6.473408e-01*S11+8.618140e+02*S12+(-1.937053e-01)*S13+4.761350e+02*S14+7.017969e-01*S15+6.890281e+00*S16+8.521027e+01*S17+(-4.849710e+01)*S18+(-1.536045e+00)*S19'
.param V38_part3='V38_part2+1.517027e+00*S20+6.012587e+01*S21+2.510038e+03*S22+1.000000e+04*S23+1.431607e+00*S24+1.000000e+04*S25+1.000000e+04*S26+1.000000e+04*S27+1.000000e+04*S28+6.608225e+02*S29'
.param V38_part4='V38_part3+(-1.689507e+01)*S30+6.484822e+01*S31+5.701237e+01*S32+2.250403e+00*S33+(-4.359748e+02)*S34+3.824810e+01*S35+1.000000e+04*S36+8.370320e+03*S37+1.000000e+04*S38+6.878651e+01*S39'
.param V38='V38_part4+(-3.400606e+00)*S40+5.877108e+01*S41+1.064799e+02*S42+1.208162e+03*S43+(-3.183862e+02)*S44'
.param V39_part1='(-6.946254e-01)*S0+8.955032e+00*S1+1.045761e+01*S2+2.242675e+00*S3+8.395883e-01*S4+2.266250e+00*S5+1.853054e+00*S6+1.803646e+01*S7+3.251546e-02*S8+7.918070e+00*S9'
.param V39_part2='V39_part1+1.253146e+00*S10+1.493781e+00*S11+4.101610e+01*S12+5.709466e-02*S13+2.859970e+01*S14+4.646856e+01*S15+9.242856e+00*S16+5.092772e+01*S17+5.176494e+01*S18+2.296837e+00*S19'
.param V39_part3='V39_part2+5.079974e+01*S20+1.426993e+01*S21+3.852381e+01*S22+4.213245e+01*S23+(-1.690381e+01)*S24+3.068290e+01*S25+5.242003e+01*S26+8.780851e+00*S27+3.552683e+01*S28+2.213468e+01*S29'
.param V39_part4='V39_part3+2.977875e+00*S30+1.893664e+01*S31+8.842465e-01*S32+1.337882e+01*S33+2.907864e+01*S34+1.534965e+01*S35+1.999515e+01*S36+3.337655e+01*S37+3.200682e+01*S38+1.238310e+01*S39'
.param V39='V39_part4+(-1.534700e+01)*S40+6.607683e+00*S41+1.739503e+01*S42+2.800879e+01*S43+1.207266e-01*S44'
.param V40_part1='9.861071e+00*S0+1.176563e+01*S1+3.544341e+01*S2+1.331228e+00*S3+1.283005e+01*S4+(-1.089974e+00)*S5+7.564778e+01*S6+5.075872e+01*S7+(-2.218949e-02)*S8+7.291403e+00*S9'
.param V40_part2='V40_part1+(-2.077834e-02)*S10+9.565433e-01*S11+9.925089e+01*S12+3.198874e-01*S13+7.288102e+01*S14+1.253803e+02*S15+1.526811e+01*S16+3.042080e+01*S17+1.969650e+01*S18+1.039287e+01*S19'
.param V40_part3='V40_part2+1.216179e+01*S20+1.439307e+02*S21+1.042619e+02*S22+4.183015e+01*S23+2.846659e+02*S24+7.240776e+01*S25+2.680592e+01*S26+1.783421e+02*S27+6.789145e+01*S28+9.322194e+01*S29'
.param V40_part4='V40_part3+9.035723e+01*S30+3.913870e+01*S31+1.701072e+01*S32+5.747224e+00*S33+1.058759e+02*S34+9.655098e+00*S35+6.800886e+01*S36+7.106179e+01*S37+8.373131e+01*S38+5.115084e+01*S39'
.param V40='V40_part4+(-9.696153e-02)*S40+(-9.043943e-01)*S41+5.150607e+01*S42+1.014980e+02*S43+1.506279e+02*S44'
.param V41_part1='(-2.139834e+00)*S0+(-6.000564e+00)*S1+(-2.499931e+01)*S2+(-2.017879e+00)*S3+(-9.791709e+00)*S4+5.172195e-01*S5+(-1.164821e+01)*S6+(-1.472217e+01)*S7+5.960495e-02*S8+(-5.049214e+00)*S9'
.param V41_part2='V41_part1+(-1.338213e+00)*S10+(-1.414177e+00)*S11+(-6.615329e+01)*S12+1.401060e-01*S13+(-8.868444e+01)*S14+(-9.018720e+01)*S15+(-7.756715e+00)*S16+(-5.714082e+01)*S17+(-3.969377e+01)*S18+(-9.934618e+00)*S19'
.param V41_part3='V41_part2+(-3.794374e+01)*S20+(-5.186064e+01)*S21+(-1.067018e+02)*S22+(-8.289679e+01)*S23+(-6.756931e+01)*S24+(-7.168924e+01)*S25+(-7.935298e+01)*S26+(-4.765156e+01)*S27+(-8.342880e+01)*S28+(-1.072433e+02)*S29'
.param V41_part4='V41_part3+(-1.532503e+01)*S30+(-4.515375e+01)*S31+(-1.322878e+01)*S32+(-1.423597e+01)*S33+(-9.411635e+01)*S34+(-2.956821e+01)*S35+(-4.056826e+01)*S36+(-7.673836e+01)*S37+(-1.077429e+02)*S38+(-2.582355e+01)*S39'
.param V41='V41_part4+7.769464e+01*S40+(-1.030486e+01)*S41+(-3.447243e+01)*S42+(-8.787128e+01)*S43+(-1.273218e+02)*S44'
.param V42_part1='1.095014e+02*S0+(-2.836868e+01)*S1+7.199703e+01*S2+(-1.231232e+02)*S3+1.959477e+02*S4+(-3.479736e+01)*S5+(-1.493834e+01)*S6+0.000000e+00*S7+0.000000e+00*S8+4.234441e+00*S9'
.param V42_part2='V42_part1+(-2.215688e+02)*S10+2.541578e+02*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+1.599405e+01*S16+0.000000e+00*S17+0.000000e+00*S18+2.391580e+02*S19'
.param V42_part3='V42_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V42_part4='V42_part3+5.339002e+01*S30+4.793884e+01*S31+1.271541e+02*S32+0.000000e+00*S33+0.000000e+00*S34+(-5.439003e+02)*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+(-4.895941e+01)*S39'
.param V42='V42_part4+1.044072e+02*S40+(-2.683863e+03)*S41+(-4.451803e+01)*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V43_part1='(-1.483303e+01)*S0+9.232443e+01*S1+(-2.211385e+01)*S2+2.029963e+02*S3+(-1.041125e+02)*S4+2.089009e+02*S5+1.000950e+02*S6+0.000000e+00*S7+0.000000e+00*S8+(-3.890025e+00)*S9'
.param V43_part2='V43_part1+1.706205e+02*S10+(-1.161013e+02)*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+(-3.902306e+01)*S16+0.000000e+00*S17+0.000000e+00*S18+(-1.907489e+02)*S19'
.param V43_part3='V43_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V43_part4='V43_part3+(-4.613226e+01)*S30+(-9.625479e+01)*S31+(-1.754460e+02)*S32+0.000000e+00*S33+0.000000e+00*S34+6.193063e+02*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+1.550525e+02*S39'
.param V43='V43_part4+3.568337e+02*S40+3.015452e+03*S41+1.008323e+02*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V44_part1='1.833209e+01*S0+3.924314e+01*S1+(-3.694009e+01)*S2+2.415398e+02*S3+(-2.773199e+01)*S4+(-8.426370e+01)*S5+9.870802e+00*S6+0.000000e+00*S7+0.000000e+00*S8+5.830383e+01*S9'
.param V44_part2='V44_part1+5.738394e+02*S10+2.211482e+01*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+4.002964e+01*S16+0.000000e+00*S17+0.000000e+00*S18+1.972591e-01*S19'
.param V44_part3='V44_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V44_part4='V44_part3+(-6.427210e+01)*S30+1.682992e+02*S31+5.609497e+02*S32+0.000000e+00*S33+0.000000e+00*S34+5.184348e+02*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+1.351412e+02*S39'
.param V44='V44_part4+(-4.750665e+02)*S40+2.882954e+03*S41+1.549971e+02*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V45_part1='0.000000e+00*S0+(-1.190045e-01)*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+(-4.729048e+00)*S5+0.000000e+00*S6+(-6.667042e-01)*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V45_part2='V45_part1+1.097388e+03*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+(-6.899878e+00)*S14+(-7.242564e-01)*S15+(-4.121888e+00)*S16+(-3.056449e+00)*S17+(-6.195416e+00)*S18+0.000000e+00*S19'
.param V45_part3='V45_part2+(-9.627185e+00)*S20+0.000000e+00*S21+0.000000e+00*S22+(-9.010603e+00)*S23+(-9.024933e-01)*S24+(-3.923694e+00)*S25+(-7.476611e+00)*S26+(-2.241656e+00)*S27+(-7.087950e+00)*S28+(-1.106303e+01)*S29'
.param V45_part4='V45_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+(-4.338511e+00)*S33+0.000000e+00*S34+0.000000e+00*S35+(-3.173155e+00)*S36+(-8.059668e+00)*S37+(-1.198917e+01)*S38+0.000000e+00*S39'
.param V45='V45_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+(-1.354909e+01)*S44'
.param V46_part1='0.000000e+00*S0+5.969654e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+2.864282e+00*S5+0.000000e+00*S6+6.782046e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V46_part2='V46_part1+1.214265e+03*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+1.365169e+01*S14+7.790900e+00*S15+3.286940e+01*S16+1.060063e+01*S17+1.633321e+01*S18+0.000000e+00*S19'
.param V46_part3='V46_part2+1.346404e+01*S20+0.000000e+00*S21+0.000000e+00*S22+1.615808e+01*S23+1.057687e+01*S24+1.308156e+01*S25+1.436377e+01*S26+1.488933e+01*S27+1.822047e+01*S28+1.854267e+01*S29'
.param V46_part4='V46_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+1.894925e+01*S33+0.000000e+00*S34+0.000000e+00*S35+1.544939e+01*S36+1.993162e+01*S37+1.929627e+01*S38+0.000000e+00*S39'
.param V46='V46_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+2.258710e+01*S44'
.param V47_part1='0.000000e+00*S0+(-3.496600e-01)*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+1.807889e+01*S5+0.000000e+00*S6+2.810494e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V47_part2='V47_part1+1.478120e+03*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+1.502558e+01*S14+2.654793e+00*S15+(-3.099553e+00)*S16+6.234852e+00*S17+1.054675e+01*S18+0.000000e+00*S19'
.param V47_part3='V47_part2+1.883507e+01*S20+0.000000e+00*S21+0.000000e+00*S22+2.273623e+01*S23+3.482932e+00*S24+1.018913e+01*S25+1.815585e+01*S26+1.018013e+01*S27+2.036060e+01*S28+3.094101e+01*S29'
.param V47_part4='V47_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+1.389242e+01*S33+0.000000e+00*S34+0.000000e+00*S35+1.399090e+01*S36+2.386769e+01*S37+3.615287e+01*S38+0.000000e+00*S39'
.param V47='V47_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+4.074264e+01*S44'
.param V48_part1='1.751227e+02*S0+4.104876e+00*S1+0.000000e+00*S2+7.330982e+02*S3+1.186421e+02*S4+4.466074e+00*S5+1.000000e+04*S6+0.000000e+00*S7+0.000000e+00*S8+3.646817e+01*S9'
.param V48_part2='V48_part1+3.462740e+03*S10+2.755434e+02*S11+5.067825e+00*S12+1.269436e+03*S13+6.905006e-01*S14+0.000000e+00*S15+1.623821e+01*S16+3.845437e-01*S17+2.281009e+00*S18+0.000000e+00*S19'
.param V48_part3='V48_part2+2.094524e+00*S20+0.000000e+00*S21+0.000000e+00*S22+1.044477e+00*S23+0.000000e+00*S24+0.000000e+00*S25+8.341777e-01*S26+1.381326e+01*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V48_part4='V48_part3+0.000000e+00*S30+3.776931e+02*S31+0.000000e+00*S32+1.863949e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+8.814833e-01*S37+8.183522e-01*S38+0.000000e+00*S39'
.param V48='V48_part4+0.000000e+00*S40+4.400800e+03*S41+6.573052e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V49_part1='3.625132e+00*S0+(-1.742596e+00)*S1+0.000000e+00*S2+7.045308e+02*S3+2.117777e+01*S4+(-1.886539e+00)*S5+(-1.000000e+04)*S6+0.000000e+00*S7+0.000000e+00*S8+2.642550e+00*S9'
.param V49_part2='V49_part1+1.830009e+02*S10+1.456208e+01*S11+(-6.920501e+00)*S12+1.269436e+03*S13+6.605727e-02*S14+0.000000e+00*S15+(-1.614170e+01)*S16+6.173023e-01*S17+(-1.834266e+00)*S18+0.000000e+00*S19'
.param V49_part3='V49_part2+(-1.437895e+00)*S20+0.000000e+00*S21+0.000000e+00*S22+(-1.747516e-01)*S23+0.000000e+00*S24+0.000000e+00*S25+(-2.761372e-01)*S26+4.221699e+01*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V49_part4='V49_part3+0.000000e+00*S30+1.280924e+02*S31+0.000000e+00*S32+(-7.830894e-01)*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+2.017903e-01*S37+(-5.504216e-02)*S38+0.000000e+00*S39'
.param V49='V49_part4+0.000000e+00*S40+1.409068e+02*S41+1.129671e+01*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V50_part1='4.102211e+01*S0+4.414808e+00*S1+0.000000e+00*S2+4.753054e+02*S3+1.029347e+01*S4+(-9.349997e-01)*S5+1.000000e+04*S6+0.000000e+00*S7+0.000000e+00*S8+3.069510e+00*S9'
.param V50_part2='V50_part1+4.427824e+02*S10+3.523387e+01*S11+(-1.822061e+00)*S12+1.269436e+03*S13+(-2.004587e-01)*S14+0.000000e+00*S15+(-6.005867e+00)*S16+(-4.312637e-01)*S17+(-1.634820e-01)*S18+0.000000e+00*S19'
.param V50_part3='V50_part2+8.795494e-02*S20+0.000000e+00*S21+0.000000e+00*S22+(-8.016884e-01)*S23+0.000000e+00*S24+0.000000e+00*S25+(-1.720932e-01)*S26+8.777617e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V50_part4='V50_part3+0.000000e+00*S30+2.556925e+02*S31+0.000000e+00*S32+6.290013e-01*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+(-1.007990e+00)*S37+(-6.493174e-01)*S38+0.000000e+00*S39'
.param V50='V50_part4+0.000000e+00*S40+1.000000e+04*S41+1.116894e+02*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V51_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+2.763392e+01*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V51_part2='V51_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+1.000000e+04*S13+0.000000e+00*S14+0.000000e+00*S15+(-6.704243e+00)*S16+0.000000e+00*S17+2.891790e+01*S18+0.000000e+00*S19'
.param V51_part3='V51_part2+(-7.116677e+00)*S20+1.000000e+04*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+6.250000e+02*S25+0.000000e+00*S26+1.000000e+04*S27+0.000000e+00*S28+2.425478e+02*S29'
.param V51_part4='V51_part3+5.888387e+03*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-9.567393e+00)*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V51='V51_part4+1.000000e+04*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+2.167352e+03*S44'
.param V52_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+(-3.208449e+01)*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V52_part2='V52_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+1.000000e+04*S13+0.000000e+00*S14+0.000000e+00*S15+1.471446e+02*S16+0.000000e+00*S17+1.359852e+02*S18+0.000000e+00*S19'
.param V52_part3='V52_part2+1.248184e+02*S20+1.000000e+04*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+6.250000e+02*S25+0.000000e+00*S26+1.000000e+04*S27+0.000000e+00*S28+1.090308e+03*S29'
.param V52_part4='V52_part3+(-7.053017e+03)*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+6.250000e+02*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V52='V52_part4+1.000000e+04*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+(-2.677884e+02)*S44'
.param V53_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+5.925499e+01*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V53_part2='V53_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+8.492323e+03*S13+0.000000e+00*S14+0.000000e+00*S15+(-3.308620e+01)*S16+0.000000e+00*S17+3.811399e+01*S18+0.000000e+00*S19'
.param V53_part3='V53_part2+8.178430e+01*S20+1.000000e+04*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+6.250000e+02*S25+0.000000e+00*S26+1.000000e+04*S27+0.000000e+00*S28+1.416876e+02*S29'
.param V53_part4='V53_part3+(-4.782898e+03)*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+5.755806e+03*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V53='V53_part4+(-1.000000e+04)*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+(-2.677884e+02)*S44'
.param _P0='V0+V1*radius_+V2*w_'
.param _P1='0.5*(_P0+sqrt(_P0*_P0+0.001))'
.param _P2='1e-09*_P1'
.param _P3='1e-09*_P1'
.param _P4='V3+V4*radius_+V5/w_'
.param _P5='0.5*(_P4+sqrt(_P4*_P4+0.001))'
.param _P6='V6+V7*radius_+V8*w_'
.param _P7='0.5*(_P6+sqrt(_P6*_P6+0.001))'
.param _P8='1e-09*_P7'
.param _P9='V9+V10*radius_+V11/w_'
.param _P10='0.5*(_P9+sqrt(_P9*_P9+0.001))'
.param _P11='V12+V13*radius_+V14*w_'
.param _P12='0.5*(_P11+sqrt(_P11*_P11+0.001))'
.param _P13='1e-09*_P12'
.param _P14='1e-09*_P12'
.param _P15='V15+V16*radius_+V17/w_'
.param _P16='0.5*(_P15+sqrt(_P15*_P15+0.001))'
.param _P17='V18+V19*radius_+V20*w_'
.param _P18='0.5*(_P17+sqrt(_P17*_P17+0.001))'
.param _P19='1e-09*_P18'
.param _P20='V21+V22*radius_+V23/w_'
.param _P21='0.5*(_P20+sqrt(_P20*_P20+0.001))'
.param _P22='V24+V25*radius_+V26*w_'
.param _P23='atan(_P22-0.5)/1.5708'
.param _P24='V27+V28*radius_+V29*w_'
.param _P25='atan(_P24-0.5)/1.5708'
.param _P26='0.5*_P23+0.5*_P25'
.param _P27='0.5*_P23-0.5*_P25'
.param _P28='V30+V31*radius_+V32*w_'
.param _P29='0.5*(_P28+sqrt(_P28*_P28+0.001))'
.param _P30='1e-15*_P29'
.param _P31='V33+V34*radius_+V35*w_'
.param _P32='0.5*(_P31+sqrt(_P31*_P31+0.001))'
.param _P33='1e-15*_P32'
.param _P34='1e-15*_P32'
.param _P35='V36+V37*radius_+V38*w_'
.param _P36='0.5*(_P35+sqrt(_P35*_P35+0.001))'
.param _P37='V39+V40*radius_+V41*w_'
.param _P38='0.5*(_P37+sqrt(_P37*_P37+0.001))'
.param _P39='V42+V43*radius_+V44*w_'
.param _P40='0.5*(_P39+sqrt(_P39*_P39+0.001))'
.param _P41='V45+V46*radius_+V47*w_'
.param _P42='0.5*(_P41+sqrt(_P41*_P41+0.001))'
.param _P43='V48+V49*radius_+V50*w_'
.param _P44='0.5*(_P43+sqrt(_P43*_P43+0.001))'
.param _P45='V51+V52*radius_+V53*w_'
.param _P46='0.5*(_P45+sqrt(_P45*_P45+0.001))'
.param _P47='1e-14*_P36'
.param _P48='100*_P38'
.param _P49='1e-15*_P40'
.param _P50='1e-14*_P36'
.param _P51='100*_P38'
.param _P52='1e-15*_P40'
.param _P53='1e-14*_P42'
.param _P54='100*_P44'
.param _P55='1e-15*_P46'
l1_sect1 PLUS _n1i_sect1 '_P2*(1+dls_3Tdiff_psub)'
l2_sect1 _n2i_sect1 MINUS '_P3*(1+dls_3Tdiff_psub)'
r1_sect1 _n1i_sect1 _n_sect1 '_P5*(1+drs_3Tdiff_psub)' tc1=0.003
r2_sect1 _n_sect1 _n2i_sect1 '_P5*(1+drs_3Tdiff_psub)' tc1=0.003
lc_sect1 _nc_sect1 CT '_P8*(1+dls_3Tdiff_psub)'
rc_sect1 _n_sect1 _nc_sect1 '_P10*(1+drs_3Tdiff_psub)' tc1=0.003
l1_sect2 PLUS _n1i_sect2 '_P13*(1+dls_3Tdiff_psub)'
l2_sect2 _n2i_sect2 MINUS '_P14*(1+dls_3Tdiff_psub)'
r1_sect2 _n1i_sect2 _n_sect2 '_P16*(1+drs_3Tdiff_psub)' tc1=0.003
r2_sect2 _n_sect2 _n2i_sect2 '_P16*(1+drs_3Tdiff_psub)' tc1=0.003
lc_sect2 _nc_sect2 CT '_P19*(1+dls_3Tdiff_psub)'
rc_sect2 _n_sect2 _nc_sect2 '_P21*(1+drs_3Tdiff_psub)' tc1=0.003
k12_sect1 l1_sect1 l2_sect1 K=_P26
k12_sect2 l1_sect2 l2_sect2 K=_P26
ks1s2_1 l1_sect1 l1_sect2 K=_P27
ks1s2_2 l2_sect1 l2_sect2 K=_P27
c12 PLUS MINUS '_P30'
c13 PLUS CT '_P33'
c23 MINUS CT '_P34'
c_1_sub PLUS _n1_1_sub '_P47'
rs_1_sub _n1_1_sub PSUB '_P48'
cs_1_sub _n1_1_sub PSUB '_P49'
c_2_sub MINUS _n1_2_sub '_P50'
rs_2_sub _n1_2_sub PSUB '_P51'
cs_2_sub _n1_2_sub PSUB '_P52'
c_3_sub CT _n1_3_sub '_P53'
rs_3_sub _n1_3_sub PSUB '_P54'
cs_3_sub _n1_3_sub PSUB '_P55'
kzero1 l1_sect1 l2_sect2 K=1e-6
kzero2 l1_sect2 l2_sect1 K=1e-6
.ends diff_ind_3t_rf_psub
