************************************************************************
* auCdl Netlist:
* 
* Library Name:  SRAM_ChargePulsation
* Top Cell Name: SRAM_CIM
* View Name:     schematic
* Netlisted on:  Jul 13 11:42:44 2022
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

.lib '/home/wangwk/projects/project_2/models_55nm/hspice/l0055ll_v1p15.lib' tt
.lib '/home/wangwk/projects/project_2/models_55nm/hspice/l0055ll_v1p15.lib' res_tt
.lib '/home/wangwk/projects/project_2/models_55nm/hspice/l0055ll_v1p15.lib' mom_tt
.options MACMOD=1

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    cell_SRAM
* View Name:    schematic
************************************************************************

.SUBCKT cell_SRAM BL Q QN SL VDD VSS WL
*.PININFO WL:I Q:O QN:O BL:B SL:B VDD:B VSS:B
XPM0 QN Q VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM1 Q QN VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XNM5 Q QN VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM4 QN Q VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM3 Q WL SL VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM2 BL WL QN VSS n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    cell_PIM
* View Name:    schematic
************************************************************************

.SUBCKT cell_PIM bl cbl in1 in2 sl vdd vss wl
*.PININFO bl:I in1:I in2:I sl:I wl:I cbl:B vdd:B vss:B
XI0 bl q qn sl vdd vss wl / cell_SRAM
XM3 net29 in1 net28 vdd p18ll_mis_ckt MR=1 L=200n W=210n
XM2 cbl in2 net29 vdd p18ll_mis_ckt MR=1 L=200n W=210n
XNM1 vdd q net28 vss n12ll_mis_ckt MR=1 L=60n W=120n
XM1 net29 qn vss vss n18ll_mis_ckt MR=1 L=200n W=210n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    cell_PIM2
* View Name:    schematic
************************************************************************

.SUBCKT cell_PIM2 bl cbl in1 in2 sl vdd vss wl
*.PININFO bl:I in1:I in2:I sl:I wl:I cbl:B vdd:B vss:B
XI0 bl q qn sl vdd vss wl / cell_SRAM
XM3 cbl in2 net9 vdd p25ll_mis_ckt MR=1 L=280n W=210n
XM2 cbl in2 net07 vdd p25ll_mis_ckt MR=1 L=280n W=210n
XM4 net9 in1 net13 vdd p25ll_mis_ckt MR=1 L=280n W=210n
XM1 net07 in1 net7 vdd p25ll_mis_ckt MR=1 L=280n W=210n
XM5 net9 qn vss vss n25ll_mis_ckt MR=1 L=280n W=210n
XM0 net07 qn vss vss n25ll_mis_ckt MR=1 L=280n W=210n
XNM3 vdd q net7 vss n12ll_mis_ckt MR=1 L=60n W=120n
XNM4 vdd q net13 vss n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    array
* View Name:    schematic
************************************************************************

.SUBCKT array bl<0> bl<1> bl<2> bl<3> bl<4> bl<5> bl<6> bl<7> bl<8> bl<9> 
+ bl<10> bl<11> bl<12> bl<13> bl<14> bl<15> bl<16> bl<17> bl<18> bl<19> bl<20> 
+ bl<21> bl<22> bl<23> bl<24> bl<25> bl<26> bl<27> bl<28> bl<29> bl<30> bl<31> 
+ bl<32> bl<33> bl<34> bl<35> bl<36> bl<37> bl<38> bl<39> bl<40> bl<41> bl<42> 
+ bl<43> bl<44> bl<45> bl<46> bl<47> bl<48> bl<49> bl<50> bl<51> bl<52> bl<53> 
+ bl<54> bl<55> bl<56> bl<57> bl<58> bl<59> bl<60> bl<61> bl<62> bl<63> 
+ blbuf<0> blbuf<1> blbuf<2> blbuf<3> blbuf<4> blbuf<5> blbuf<6> blbuf<7> 
+ blbuf<8> blbuf<9> blbuf<10> blbuf<11> blbuf<12> blbuf<13> blbuf<14> 
+ blbuf<15> cbl<0> cbl<1> cbl<2> cbl<3> cbl<4> cbl<5> cbl<6> cbl<7> cbl<8> 
+ cbl<9> cbl<10> cbl<11> cbl<12> cbl<13> cbl<14> cbl<15> cbl<16> cbl<17> 
+ cbl<18> cbl<19> cbl<20> cbl<21> cbl<22> cbl<23> cbl<24> cbl<25> cbl<26> 
+ cbl<27> cbl<28> cbl<29> cbl<30> cbl<31> in1<0> in1<1> in1<2> in1<3> in1<4> 
+ in1<5> in1<6> in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> 
+ in1<15> in1<16> in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> 
+ in1<24> in1<25> in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> 
+ in1<33> in1<34> in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> 
+ in1<42> in1<43> in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> 
+ in1<51> in1<52> in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> 
+ in1<60> in1<61> in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> 
+ in1<69> in1<70> in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> 
+ in1<78> in1<79> in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> 
+ in1<87> in1<88> in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> 
+ in1<96> in1<97> in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> 
+ in1<105> in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> 
+ in1<113> in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> 
+ in1<121> in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> 
+ in2<2> in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> 
+ in2<12> in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> 
+ in2<21> in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> 
+ in2<30> in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> 
+ in2<39> in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> 
+ in2<48> in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> 
+ in2<57> in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> 
+ in2<66> in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> 
+ in2<75> in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> 
+ in2<84> in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> 
+ in2<93> in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> 
+ in2<102> in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> 
+ in2<110> in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> 
+ in2<118> in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> 
+ in2<126> in2<127> sl<0> sl<1> sl<2> sl<3> sl<4> sl<5> sl<6> sl<7> sl<8> 
+ sl<9> sl<10> sl<11> sl<12> sl<13> sl<14> sl<15> sl<16> sl<17> sl<18> sl<19> 
+ sl<20> sl<21> sl<22> sl<23> sl<24> sl<25> sl<26> sl<27> sl<28> sl<29> sl<30> 
+ sl<31> sl<32> sl<33> sl<34> sl<35> sl<36> sl<37> sl<38> sl<39> sl<40> sl<41> 
+ sl<42> sl<43> sl<44> sl<45> sl<46> sl<47> sl<48> sl<49> sl<50> sl<51> sl<52> 
+ sl<53> sl<54> sl<55> sl<56> sl<57> sl<58> sl<59> sl<60> sl<61> sl<62> sl<63> 
+ slbuf<0> slbuf<1> slbuf<2> slbuf<3> slbuf<4> slbuf<5> slbuf<6> slbuf<7> 
+ slbuf<8> slbuf<9> slbuf<10> slbuf<11> slbuf<12> slbuf<13> slbuf<14> 
+ slbuf<15> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> 
+ wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> 
+ wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> 
+ wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> 
+ wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> 
+ wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> 
+ wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> 
+ wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> 
+ wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> 
+ wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127>
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I bl<4>:I bl<5>:I bl<6>:I bl<7>:I 
*.PININFO bl<8>:I bl<9>:I bl<10>:I bl<11>:I bl<12>:I bl<13>:I bl<14>:I 
*.PININFO bl<15>:I bl<16>:I bl<17>:I bl<18>:I bl<19>:I bl<20>:I bl<21>:I 
*.PININFO bl<22>:I bl<23>:I bl<24>:I bl<25>:I bl<26>:I bl<27>:I bl<28>:I 
*.PININFO bl<29>:I bl<30>:I bl<31>:I bl<32>:I bl<33>:I bl<34>:I bl<35>:I 
*.PININFO bl<36>:I bl<37>:I bl<38>:I bl<39>:I bl<40>:I bl<41>:I bl<42>:I 
*.PININFO bl<43>:I bl<44>:I bl<45>:I bl<46>:I bl<47>:I bl<48>:I bl<49>:I 
*.PININFO bl<50>:I bl<51>:I bl<52>:I bl<53>:I bl<54>:I bl<55>:I bl<56>:I 
*.PININFO bl<57>:I bl<58>:I bl<59>:I bl<60>:I bl<61>:I bl<62>:I bl<63>:I 
*.PININFO in1<0>:I in1<1>:I in1<2>:I in1<3>:I in1<4>:I in1<5>:I in1<6>:I 
*.PININFO in1<7>:I in1<8>:I in1<9>:I in1<10>:I in1<11>:I in1<12>:I in1<13>:I 
*.PININFO in1<14>:I in1<15>:I in1<16>:I in1<17>:I in1<18>:I in1<19>:I 
*.PININFO in1<20>:I in1<21>:I in1<22>:I in1<23>:I in1<24>:I in1<25>:I 
*.PININFO in1<26>:I in1<27>:I in1<28>:I in1<29>:I in1<30>:I in1<31>:I 
*.PININFO in1<32>:I in1<33>:I in1<34>:I in1<35>:I in1<36>:I in1<37>:I 
*.PININFO in1<38>:I in1<39>:I in1<40>:I in1<41>:I in1<42>:I in1<43>:I 
*.PININFO in1<44>:I in1<45>:I in1<46>:I in1<47>:I in1<48>:I in1<49>:I 
*.PININFO in1<50>:I in1<51>:I in1<52>:I in1<53>:I in1<54>:I in1<55>:I 
*.PININFO in1<56>:I in1<57>:I in1<58>:I in1<59>:I in1<60>:I in1<61>:I 
*.PININFO in1<62>:I in1<63>:I in1<64>:I in1<65>:I in1<66>:I in1<67>:I 
*.PININFO in1<68>:I in1<69>:I in1<70>:I in1<71>:I in1<72>:I in1<73>:I 
*.PININFO in1<74>:I in1<75>:I in1<76>:I in1<77>:I in1<78>:I in1<79>:I 
*.PININFO in1<80>:I in1<81>:I in1<82>:I in1<83>:I in1<84>:I in1<85>:I 
*.PININFO in1<86>:I in1<87>:I in1<88>:I in1<89>:I in1<90>:I in1<91>:I 
*.PININFO in1<92>:I in1<93>:I in1<94>:I in1<95>:I in1<96>:I in1<97>:I 
*.PININFO in1<98>:I in1<99>:I in1<100>:I in1<101>:I in1<102>:I in1<103>:I 
*.PININFO in1<104>:I in1<105>:I in1<106>:I in1<107>:I in1<108>:I in1<109>:I 
*.PININFO in1<110>:I in1<111>:I in1<112>:I in1<113>:I in1<114>:I in1<115>:I 
*.PININFO in1<116>:I in1<117>:I in1<118>:I in1<119>:I in1<120>:I in1<121>:I 
*.PININFO in1<122>:I in1<123>:I in1<124>:I in1<125>:I in1<126>:I in1<127>:I 
*.PININFO in2<0>:I in2<1>:I in2<2>:I in2<3>:I in2<4>:I in2<5>:I in2<6>:I 
*.PININFO in2<7>:I in2<8>:I in2<9>:I in2<10>:I in2<11>:I in2<12>:I in2<13>:I 
*.PININFO in2<14>:I in2<15>:I in2<16>:I in2<17>:I in2<18>:I in2<19>:I 
*.PININFO in2<20>:I in2<21>:I in2<22>:I in2<23>:I in2<24>:I in2<25>:I 
*.PININFO in2<26>:I in2<27>:I in2<28>:I in2<29>:I in2<30>:I in2<31>:I 
*.PININFO in2<32>:I in2<33>:I in2<34>:I in2<35>:I in2<36>:I in2<37>:I 
*.PININFO in2<38>:I in2<39>:I in2<40>:I in2<41>:I in2<42>:I in2<43>:I 
*.PININFO in2<44>:I in2<45>:I in2<46>:I in2<47>:I in2<48>:I in2<49>:I 
*.PININFO in2<50>:I in2<51>:I in2<52>:I in2<53>:I in2<54>:I in2<55>:I 
*.PININFO in2<56>:I in2<57>:I in2<58>:I in2<59>:I in2<60>:I in2<61>:I 
*.PININFO in2<62>:I in2<63>:I in2<64>:I in2<65>:I in2<66>:I in2<67>:I 
*.PININFO in2<68>:I in2<69>:I in2<70>:I in2<71>:I in2<72>:I in2<73>:I 
*.PININFO in2<74>:I in2<75>:I in2<76>:I in2<77>:I in2<78>:I in2<79>:I 
*.PININFO in2<80>:I in2<81>:I in2<82>:I in2<83>:I in2<84>:I in2<85>:I 
*.PININFO in2<86>:I in2<87>:I in2<88>:I in2<89>:I in2<90>:I in2<91>:I 
*.PININFO in2<92>:I in2<93>:I in2<94>:I in2<95>:I in2<96>:I in2<97>:I 
*.PININFO in2<98>:I in2<99>:I in2<100>:I in2<101>:I in2<102>:I in2<103>:I 
*.PININFO in2<104>:I in2<105>:I in2<106>:I in2<107>:I in2<108>:I in2<109>:I 
*.PININFO in2<110>:I in2<111>:I in2<112>:I in2<113>:I in2<114>:I in2<115>:I 
*.PININFO in2<116>:I in2<117>:I in2<118>:I in2<119>:I in2<120>:I in2<121>:I 
*.PININFO in2<122>:I in2<123>:I in2<124>:I in2<125>:I in2<126>:I in2<127>:I 
*.PININFO sl<0>:I sl<1>:I sl<2>:I sl<3>:I sl<4>:I sl<5>:I sl<6>:I sl<7>:I 
*.PININFO sl<8>:I sl<9>:I sl<10>:I sl<11>:I sl<12>:I sl<13>:I sl<14>:I 
*.PININFO sl<15>:I sl<16>:I sl<17>:I sl<18>:I sl<19>:I sl<20>:I sl<21>:I 
*.PININFO sl<22>:I sl<23>:I sl<24>:I sl<25>:I sl<26>:I sl<27>:I sl<28>:I 
*.PININFO sl<29>:I sl<30>:I sl<31>:I sl<32>:I sl<33>:I sl<34>:I sl<35>:I 
*.PININFO sl<36>:I sl<37>:I sl<38>:I sl<39>:I sl<40>:I sl<41>:I sl<42>:I 
*.PININFO sl<43>:I sl<44>:I sl<45>:I sl<46>:I sl<47>:I sl<48>:I sl<49>:I 
*.PININFO sl<50>:I sl<51>:I sl<52>:I sl<53>:I sl<54>:I sl<55>:I sl<56>:I 
*.PININFO sl<57>:I sl<58>:I sl<59>:I sl<60>:I sl<61>:I sl<62>:I sl<63>:I 
*.PININFO wl<0>:I wl<1>:I wl<2>:I wl<3>:I wl<4>:I wl<5>:I wl<6>:I wl<7>:I 
*.PININFO wl<8>:I wl<9>:I wl<10>:I wl<11>:I wl<12>:I wl<13>:I wl<14>:I 
*.PININFO wl<15>:I wl<16>:I wl<17>:I wl<18>:I wl<19>:I wl<20>:I wl<21>:I 
*.PININFO wl<22>:I wl<23>:I wl<24>:I wl<25>:I wl<26>:I wl<27>:I wl<28>:I 
*.PININFO wl<29>:I wl<30>:I wl<31>:I wl<32>:I wl<33>:I wl<34>:I wl<35>:I 
*.PININFO wl<36>:I wl<37>:I wl<38>:I wl<39>:I wl<40>:I wl<41>:I wl<42>:I 
*.PININFO wl<43>:I wl<44>:I wl<45>:I wl<46>:I wl<47>:I wl<48>:I wl<49>:I 
*.PININFO wl<50>:I wl<51>:I wl<52>:I wl<53>:I wl<54>:I wl<55>:I wl<56>:I 
*.PININFO wl<57>:I wl<58>:I wl<59>:I wl<60>:I wl<61>:I wl<62>:I wl<63>:I 
*.PININFO wl<64>:I wl<65>:I wl<66>:I wl<67>:I wl<68>:I wl<69>:I wl<70>:I 
*.PININFO wl<71>:I wl<72>:I wl<73>:I wl<74>:I wl<75>:I wl<76>:I wl<77>:I 
*.PININFO wl<78>:I wl<79>:I wl<80>:I wl<81>:I wl<82>:I wl<83>:I wl<84>:I 
*.PININFO wl<85>:I wl<86>:I wl<87>:I wl<88>:I wl<89>:I wl<90>:I wl<91>:I 
*.PININFO wl<92>:I wl<93>:I wl<94>:I wl<95>:I wl<96>:I wl<97>:I wl<98>:I 
*.PININFO wl<99>:I wl<100>:I wl<101>:I wl<102>:I wl<103>:I wl<104>:I wl<105>:I 
*.PININFO wl<106>:I wl<107>:I wl<108>:I wl<109>:I wl<110>:I wl<111>:I 
*.PININFO wl<112>:I wl<113>:I wl<114>:I wl<115>:I wl<116>:I wl<117>:I 
*.PININFO wl<118>:I wl<119>:I wl<120>:I wl<121>:I wl<122>:I wl<123>:I 
*.PININFO wl<124>:I wl<125>:I wl<126>:I wl<127>:I blbuf<0>:B blbuf<1>:B 
*.PININFO blbuf<2>:B blbuf<3>:B blbuf<4>:B blbuf<5>:B blbuf<6>:B blbuf<7>:B 
*.PININFO blbuf<8>:B blbuf<9>:B blbuf<10>:B blbuf<11>:B blbuf<12>:B 
*.PININFO blbuf<13>:B blbuf<14>:B blbuf<15>:B cbl<0>:B cbl<1>:B cbl<2>:B 
*.PININFO cbl<3>:B cbl<4>:B cbl<5>:B cbl<6>:B cbl<7>:B cbl<8>:B cbl<9>:B 
*.PININFO cbl<10>:B cbl<11>:B cbl<12>:B cbl<13>:B cbl<14>:B cbl<15>:B 
*.PININFO cbl<16>:B cbl<17>:B cbl<18>:B cbl<19>:B cbl<20>:B cbl<21>:B 
*.PININFO cbl<22>:B cbl<23>:B cbl<24>:B cbl<25>:B cbl<26>:B cbl<27>:B 
*.PININFO cbl<28>:B cbl<29>:B cbl<30>:B cbl<31>:B slbuf<0>:B slbuf<1>:B 
*.PININFO slbuf<2>:B slbuf<3>:B slbuf<4>:B slbuf<5>:B slbuf<6>:B slbuf<7>:B 
*.PININFO slbuf<8>:B slbuf<9>:B slbuf<10>:B slbuf<11>:B slbuf<12>:B 
*.PININFO slbuf<13>:B slbuf<14>:B slbuf<15>:B vdd:B vss:B
XI17168 bl<2> cbl<1> in1<61> in2<61> sl<2> vdd vss wl<61> / cell_PIM
XI17166 bl<2> cbl<1> in1<59> in2<59> sl<2> vdd vss wl<59> / cell_PIM
XI17167 bl<2> cbl<1> in1<60> in2<60> sl<2> vdd vss wl<60> / cell_PIM
XI25357 vss vss in1<0> in2<0> vss vdd vss wl<0> / cell_PIM
XI25358 vss vss vdd vdd vss vdd vss vss / cell_PIM
XI25354 vss vss in1<4> in2<4> vss vdd vss wl<4> / cell_PIM
XI25355 vss vss in1<1> in2<1> vss vdd vss wl<1> / cell_PIM
XI25356 vss vss in1<2> in2<2> vss vdd vss wl<2> / cell_PIM
XI24707 bl<62> cbl<31> in1<11> in2<11> sl<62> vdd vss wl<11> / cell_PIM
XI24708 bl<62> cbl<31> in1<9> in2<9> sl<62> vdd vss wl<9> / cell_PIM
XI24705 bl<62> cbl<31> in1<10> in2<10> sl<62> vdd vss wl<10> / cell_PIM
XI24706 bl<62> cbl<31> in1<12> in2<12> sl<62> vdd vss wl<12> / cell_PIM
XI24057 bl<54> cbl<27> in1<29> in2<29> sl<54> vdd vss wl<29> / cell_PIM
XI24058 bl<54> cbl<27> in1<31> in2<31> sl<54> vdd vss wl<31> / cell_PIM
XI22884 bl<62> cbl<31> in1<66> in2<66> sl<62> vdd vss wl<66> / cell_PIM
XI22885 bl<62> cbl<31> in1<65> in2<65> sl<62> vdd vss wl<65> / cell_PIM
XI22237 bl<54> cbl<27> in1<84> in2<84> sl<54> vdd vss wl<84> / cell_PIM
XI22234 bl<54> cbl<27> in1<88> in2<88> sl<54> vdd vss wl<88> / cell_PIM
XI22235 bl<54> cbl<27> in1<86> in2<86> sl<54> vdd vss wl<86> / cell_PIM
XI22236 bl<54> cbl<27> in1<85> in2<85> sl<54> vdd vss wl<85> / cell_PIM
XI21587 bl<50> cbl<25> in1<106> in2<106> sl<50> vdd vss wl<106> / cell_PIM
XI21588 bl<50> cbl<25> in1<107> in2<107> sl<50> vdd vss wl<107> / cell_PIM
XI20937 bl<44> cbl<22> in1<125> in2<125> sl<44> vdd vss wl<125> / cell_PIM
XI20938 bl<44> cbl<22> in1<126> in2<126> sl<44> vdd vss wl<126> / cell_PIM
XI20935 bl<44> cbl<22> in1<123> in2<123> sl<44> vdd vss wl<123> / cell_PIM
XI20936 bl<44> cbl<22> in1<124> in2<124> sl<44> vdd vss wl<124> / cell_PIM
XI20285 bl<16> cbl<8> in1<36> in2<36> sl<16> vdd vss wl<36> / cell_PIM
XI20286 bl<16> cbl<8> in1<32> in2<32> sl<16> vdd vss wl<32> / cell_PIM
XI20287 bl<16> cbl<8> in1<33> in2<33> sl<16> vdd vss wl<33> / cell_PIM
XI19767 bl<18> cbl<9> in1<67> in2<67> sl<18> vdd vss wl<67> / cell_PIM
XI19768 bl<18> cbl<9> in1<66> in2<66> sl<18> vdd vss wl<66> / cell_PIM
XI19765 bl<18> cbl<9> in1<68> in2<68> sl<18> vdd vss wl<68> / cell_PIM
XI19766 bl<18> cbl<9> in1<69> in2<69> sl<18> vdd vss wl<69> / cell_PIM
XI19117 bl<26> cbl<13> in1<111> in2<111> sl<26> vdd vss wl<111> / cell_PIM
XI19118 bl<26> cbl<13> in1<112> in2<112> sl<26> vdd vss wl<112> / cell_PIM
XI18467 bl<14> cbl<7> in1<44> in2<44> sl<14> vdd vss wl<44> / cell_PIM
XI18468 bl<14> cbl<7> in1<47> in2<47> sl<14> vdd vss wl<47> / cell_PIM
XI17817 bl<12> cbl<6> in1<127> in2<127> sl<12> vdd vss wl<127> / cell_PIM
XI17815 bl<12> cbl<6> in1<125> in2<125> sl<12> vdd vss wl<125> / cell_PIM
XI17816 bl<12> cbl<6> in1<126> in2<126> sl<12> vdd vss wl<126> / cell_PIM
XI16821 bl<0> cbl<0> in1<42> in2<42> sl<0> vdd vss wl<42> / cell_PIM
XI16822 bl<0> cbl<0> in1<43> in2<43> sl<0> vdd vss wl<43> / cell_PIM
XI16820 bl<0> cbl<0> in1<41> in2<41> sl<0> vdd vss wl<41> / cell_PIM
XI24709 bl<62> cbl<31> in1<8> in2<8> sl<62> vdd vss wl<8> / cell_PIM
XI24060 bl<54> cbl<27> in1<28> in2<28> sl<54> vdd vss wl<28> / cell_PIM
XI24061 bl<54> cbl<27> in1<27> in2<27> sl<54> vdd vss wl<27> / cell_PIM
XI24059 bl<54> cbl<27> in1<30> in2<30> sl<54> vdd vss wl<30> / cell_PIM
XI23410 bl<46> cbl<23> in1<50> in2<50> sl<46> vdd vss wl<50> / cell_PIM
XI23411 bl<46> cbl<23> in1<49> in2<49> sl<46> vdd vss wl<49> / cell_PIM
XI23412 bl<46> cbl<23> in1<47> in2<47> sl<46> vdd vss wl<47> / cell_PIM
XI23413 bl<46> cbl<23> in1<46> in2<46> sl<46> vdd vss wl<46> / cell_PIM
XI23409 bl<46> cbl<23> in1<48> in2<48> sl<46> vdd vss wl<48> / cell_PIM
XI22891 bl<32> cbl<16> in1<63> in2<63> sl<32> vdd vss wl<63> / cell_PIM
XI22892 bl<32> cbl<16> in1<64> in2<64> sl<32> vdd vss wl<64> / cell_PIM
XI22243 bl<56> cbl<28> in1<87> in2<87> sl<56> vdd vss wl<87> / cell_PIM
XI21590 bl<50> cbl<25> in1<104> in2<104> sl<50> vdd vss wl<104> / cell_PIM
XI21589 bl<50> cbl<25> in1<105> in2<105> sl<50> vdd vss wl<105> / cell_PIM
XI20939 bl<44> cbl<22> in1<127> in2<127> sl<44> vdd vss wl<127> / cell_PIM
XI20293 bl<18> cbl<9> in1<34> in2<34> sl<18> vdd vss wl<34> / cell_PIM
XI19769 bl<18> cbl<9> in1<65> in2<65> sl<18> vdd vss wl<65> / cell_PIM
XI19120 bl<26> cbl<13> in1<109> in2<109> sl<26> vdd vss wl<109> / cell_PIM
XI19121 bl<26> cbl<13> in1<108> in2<108> sl<26> vdd vss wl<108> / cell_PIM
XI19119 bl<26> cbl<13> in1<110> in2<110> sl<26> vdd vss wl<110> / cell_PIM
XI18470 bl<14> cbl<7> in1<45> in2<45> sl<14> vdd vss wl<45> / cell_PIM
XI18469 bl<14> cbl<7> in1<46> in2<46> sl<14> vdd vss wl<46> / cell_PIM
XI17821 bl<14> cbl<7> in1<125> in2<125> sl<14> vdd vss wl<125> / cell_PIM
XI17822 bl<14> cbl<7> in1<126> in2<126> sl<14> vdd vss wl<126> / cell_PIM
XI17823 bl<14> cbl<7> in1<127> in2<127> sl<14> vdd vss wl<127> / cell_PIM
XI17169 bl<2> cbl<1> in1<62> in2<62> sl<2> vdd vss wl<62> / cell_PIM
XI17165 bl<2> cbl<1> in1<58> in2<58> sl<2> vdd vss wl<58> / cell_PIM
XI17159 bl<2> cbl<1> in1<67> in2<67> sl<2> vdd vss wl<67> / cell_PIM
XI17156 bl<2> cbl<1> in1<64> in2<64> sl<2> vdd vss wl<64> / cell_PIM
XI17150 bl<2> cbl<1> in1<71> in2<71> sl<2> vdd vss wl<71> / cell_PIM
XI17147 bl<2> cbl<1> in1<68> in2<68> sl<2> vdd vss wl<68> / cell_PIM
XI17141 bl<2> cbl<1> in1<76> in2<76> sl<2> vdd vss wl<76> / cell_PIM
XI17138 bl<2> cbl<1> in1<73> in2<73> sl<2> vdd vss wl<73> / cell_PIM
XI17129 bl<2> cbl<1> in1<79> in2<79> sl<2> vdd vss wl<79> / cell_PIM
XI17120 bl<2> cbl<1> in1<85> in2<85> sl<2> vdd vss wl<85> / cell_PIM
XI17117 bl<2> cbl<1> in1<82> in2<82> sl<2> vdd vss wl<82> / cell_PIM
XI17111 bl<2> cbl<1> in1<91> in2<91> sl<2> vdd vss wl<91> / cell_PIM
XI17108 bl<2> cbl<1> in1<88> in2<88> sl<2> vdd vss wl<88> / cell_PIM
XI17102 bl<2> cbl<1> in1<95> in2<95> sl<2> vdd vss wl<95> / cell_PIM
XI17099 bl<2> cbl<1> in1<92> in2<92> sl<2> vdd vss wl<92> / cell_PIM
XI17093 bl<2> cbl<1> in1<100> in2<100> sl<2> vdd vss wl<100> / cell_PIM
XI17090 bl<2> cbl<1> in1<97> in2<97> sl<2> vdd vss wl<97> / cell_PIM
XI17081 bl<2> cbl<1> in1<103> in2<103> sl<2> vdd vss wl<103> / cell_PIM
XI17072 bl<2> cbl<1> in1<109> in2<109> sl<2> vdd vss wl<109> / cell_PIM
XI17069 bl<2> cbl<1> in1<106> in2<106> sl<2> vdd vss wl<106> / cell_PIM
XI17063 bl<2> cbl<1> in1<115> in2<115> sl<2> vdd vss wl<115> / cell_PIM
XI17060 bl<2> cbl<1> in1<112> in2<112> sl<2> vdd vss wl<112> / cell_PIM
XI17054 bl<2> cbl<1> in1<119> in2<119> sl<2> vdd vss wl<119> / cell_PIM
XI17051 bl<2> cbl<1> in1<116> in2<116> sl<2> vdd vss wl<116> / cell_PIM
XI17045 bl<2> cbl<1> in1<124> in2<124> sl<2> vdd vss wl<124> / cell_PIM
XI17042 bl<2> cbl<1> in1<121> in2<121> sl<2> vdd vss wl<121> / cell_PIM
XI17035 bl<2> cbl<1> in1<125> in2<125> sl<2> vdd vss wl<125> / cell_PIM
XI16905 bl<0> cbl<0> in1<126> in2<126> sl<0> vdd vss wl<126> / cell_PIM
XI16902 bl<0> cbl<0> in1<123> in2<123> sl<0> vdd vss wl<123> / cell_PIM
XI16899 bl<0> cbl<0> in1<120> in2<120> sl<0> vdd vss wl<120> / cell_PIM
XI16896 bl<0> cbl<0> in1<117> in2<117> sl<0> vdd vss wl<117> / cell_PIM
XI16893 bl<0> cbl<0> in1<114> in2<114> sl<0> vdd vss wl<114> / cell_PIM
XI16890 bl<0> cbl<0> in1<111> in2<111> sl<0> vdd vss wl<111> / cell_PIM
XI16887 bl<0> cbl<0> in1<108> in2<108> sl<0> vdd vss wl<108> / cell_PIM
XI16884 bl<0> cbl<0> in1<105> in2<105> sl<0> vdd vss wl<105> / cell_PIM
XI16881 bl<0> cbl<0> in1<102> in2<102> sl<0> vdd vss wl<102> / cell_PIM
XI16878 bl<0> cbl<0> in1<99> in2<99> sl<0> vdd vss wl<99> / cell_PIM
XI16875 bl<0> cbl<0> in1<96> in2<96> sl<0> vdd vss wl<96> / cell_PIM
XI16872 bl<0> cbl<0> in1<93> in2<93> sl<0> vdd vss wl<93> / cell_PIM
XI16869 bl<0> cbl<0> in1<90> in2<90> sl<0> vdd vss wl<90> / cell_PIM
XI16866 bl<0> cbl<0> in1<87> in2<87> sl<0> vdd vss wl<87> / cell_PIM
XI16863 bl<0> cbl<0> in1<84> in2<84> sl<0> vdd vss wl<84> / cell_PIM
XI16860 bl<0> cbl<0> in1<81> in2<81> sl<0> vdd vss wl<81> / cell_PIM
XI16857 bl<0> cbl<0> in1<78> in2<78> sl<0> vdd vss wl<78> / cell_PIM
XI16854 bl<0> cbl<0> in1<75> in2<75> sl<0> vdd vss wl<75> / cell_PIM
XI16851 bl<0> cbl<0> in1<72> in2<72> sl<0> vdd vss wl<72> / cell_PIM
XI16848 bl<0> cbl<0> in1<69> in2<69> sl<0> vdd vss wl<69> / cell_PIM
XI16810 bl<0> cbl<0> in1<31> in2<31> sl<0> vdd vss wl<31> / cell_PIM
XI16807 bl<0> cbl<0> in1<28> in2<28> sl<0> vdd vss wl<28> / cell_PIM
XI16804 bl<0> cbl<0> in1<25> in2<25> sl<0> vdd vss wl<25> / cell_PIM
XI16801 bl<0> cbl<0> in1<22> in2<22> sl<0> vdd vss wl<22> / cell_PIM
XI16798 bl<0> cbl<0> in1<19> in2<19> sl<0> vdd vss wl<19> / cell_PIM
XI16795 bl<0> cbl<0> in1<16> in2<16> sl<0> vdd vss wl<16> / cell_PIM
XI16792 bl<0> cbl<0> in1<13> in2<13> sl<0> vdd vss wl<13> / cell_PIM
XI16789 bl<0> cbl<0> in1<10> in2<10> sl<0> vdd vss wl<10> / cell_PIM
XI16786 bl<0> cbl<0> in1<7> in2<7> sl<0> vdd vss wl<7> / cell_PIM
XI16783 bl<0> cbl<0> in1<4> in2<4> sl<0> vdd vss wl<4> / cell_PIM
XI16780 bl<0> cbl<0> in1<1> in2<1> sl<0> vdd vss wl<1> / cell_PIM
XI16846 bl<0> cbl<0> in1<67> in2<67> sl<0> vdd vss wl<67> / cell_PIM
XI16843 bl<0> cbl<0> in1<64> in2<64> sl<0> vdd vss wl<64> / cell_PIM
XI16840 bl<0> cbl<0> in1<61> in2<61> sl<0> vdd vss wl<61> / cell_PIM
XI16837 bl<0> cbl<0> in1<58> in2<58> sl<0> vdd vss wl<58> / cell_PIM
XI16834 bl<0> cbl<0> in1<55> in2<55> sl<0> vdd vss wl<55> / cell_PIM
XI16831 bl<0> cbl<0> in1<52> in2<52> sl<0> vdd vss wl<52> / cell_PIM
XI16828 bl<0> cbl<0> in1<49> in2<49> sl<0> vdd vss wl<49> / cell_PIM
XI16825 bl<0> cbl<0> in1<46> in2<46> sl<0> vdd vss wl<46> / cell_PIM
XI16819 bl<0> cbl<0> in1<40> in2<40> sl<0> vdd vss wl<40> / cell_PIM
XI16818 bl<0> cbl<0> in1<39> in2<39> sl<0> vdd vss wl<39> / cell_PIM
XI16817 bl<0> cbl<0> in1<38> in2<38> sl<0> vdd vss wl<38> / cell_PIM
XI17158 bl<2> cbl<1> in1<66> in2<66> sl<2> vdd vss wl<66> / cell_PIM
XI17157 bl<2> cbl<1> in1<65> in2<65> sl<2> vdd vss wl<65> / cell_PIM
XI17155 bl<2> cbl<1> in1<63> in2<63> sl<2> vdd vss wl<63> / cell_PIM
XI17149 bl<2> cbl<1> in1<70> in2<70> sl<2> vdd vss wl<70> / cell_PIM
XI17148 bl<2> cbl<1> in1<69> in2<69> sl<2> vdd vss wl<69> / cell_PIM
XI17140 bl<2> cbl<1> in1<75> in2<75> sl<2> vdd vss wl<75> / cell_PIM
XI17139 bl<2> cbl<1> in1<74> in2<74> sl<2> vdd vss wl<74> / cell_PIM
XI17137 bl<2> cbl<1> in1<72> in2<72> sl<2> vdd vss wl<72> / cell_PIM
XI17131 bl<2> cbl<1> in1<81> in2<81> sl<2> vdd vss wl<81> / cell_PIM
XI17130 bl<2> cbl<1> in1<80> in2<80> sl<2> vdd vss wl<80> / cell_PIM
XI17128 bl<2> cbl<1> in1<78> in2<78> sl<2> vdd vss wl<78> / cell_PIM
XI17127 bl<2> cbl<1> in1<77> in2<77> sl<2> vdd vss wl<77> / cell_PIM
XI17121 bl<2> cbl<1> in1<86> in2<86> sl<2> vdd vss wl<86> / cell_PIM
XI17119 bl<2> cbl<1> in1<84> in2<84> sl<2> vdd vss wl<84> / cell_PIM
XI17118 bl<2> cbl<1> in1<83> in2<83> sl<2> vdd vss wl<83> / cell_PIM
XI17110 bl<2> cbl<1> in1<90> in2<90> sl<2> vdd vss wl<90> / cell_PIM
XI17109 bl<2> cbl<1> in1<89> in2<89> sl<2> vdd vss wl<89> / cell_PIM
XI17107 bl<2> cbl<1> in1<87> in2<87> sl<2> vdd vss wl<87> / cell_PIM
XI17101 bl<2> cbl<1> in1<94> in2<94> sl<2> vdd vss wl<94> / cell_PIM
XI17100 bl<2> cbl<1> in1<93> in2<93> sl<2> vdd vss wl<93> / cell_PIM
XI17092 bl<2> cbl<1> in1<99> in2<99> sl<2> vdd vss wl<99> / cell_PIM
XI17091 bl<2> cbl<1> in1<98> in2<98> sl<2> vdd vss wl<98> / cell_PIM
XI17089 bl<2> cbl<1> in1<96> in2<96> sl<2> vdd vss wl<96> / cell_PIM
XI17083 bl<2> cbl<1> in1<105> in2<105> sl<2> vdd vss wl<105> / cell_PIM
XI17082 bl<2> cbl<1> in1<104> in2<104> sl<2> vdd vss wl<104> / cell_PIM
XI17080 bl<2> cbl<1> in1<102> in2<102> sl<2> vdd vss wl<102> / cell_PIM
XI17079 bl<2> cbl<1> in1<101> in2<101> sl<2> vdd vss wl<101> / cell_PIM
XI17073 bl<2> cbl<1> in1<110> in2<110> sl<2> vdd vss wl<110> / cell_PIM
XI17071 bl<2> cbl<1> in1<108> in2<108> sl<2> vdd vss wl<108> / cell_PIM
XI17070 bl<2> cbl<1> in1<107> in2<107> sl<2> vdd vss wl<107> / cell_PIM
XI17062 bl<2> cbl<1> in1<114> in2<114> sl<2> vdd vss wl<114> / cell_PIM
XI17061 bl<2> cbl<1> in1<113> in2<113> sl<2> vdd vss wl<113> / cell_PIM
XI17059 bl<2> cbl<1> in1<111> in2<111> sl<2> vdd vss wl<111> / cell_PIM
XI17053 bl<2> cbl<1> in1<118> in2<118> sl<2> vdd vss wl<118> / cell_PIM
XI17052 bl<2> cbl<1> in1<117> in2<117> sl<2> vdd vss wl<117> / cell_PIM
XI17044 bl<2> cbl<1> in1<123> in2<123> sl<2> vdd vss wl<123> / cell_PIM
XI17043 bl<2> cbl<1> in1<122> in2<122> sl<2> vdd vss wl<122> / cell_PIM
XI17041 bl<2> cbl<1> in1<120> in2<120> sl<2> vdd vss wl<120> / cell_PIM
XI17036 bl<2> cbl<1> in1<126> in2<126> sl<2> vdd vss wl<126> / cell_PIM
XI25352 vss vss in1<7> in2<7> vss vdd vss wl<7> / cell_PIM
XI25351 vss vss in1<6> in2<6> vss vdd vss wl<6> / cell_PIM
XI25350 vss vss in1<5> in2<5> vss vdd vss wl<5> / cell_PIM
XI25349 vss vss in1<9> in2<9> vss vdd vss wl<9> / cell_PIM
XI25353 vss vss in1<3> in2<3> vss vdd vss wl<3> / cell_PIM
XI25348 vss vss in1<8> in2<8> vss vdd vss wl<8> / cell_PIM
XI25347 vss vss in1<11> in2<11> vss vdd vss wl<11> / cell_PIM
XI25346 vss vss in1<10> in2<10> vss vdd vss wl<10> / cell_PIM
XI25345 vss vss in1<12> in2<12> vss vdd vss wl<12> / cell_PIM
XI25344 vss vss in1<14> in2<14> vss vdd vss wl<14> / cell_PIM
XI24698 bl<60> cbl<30> in1<8> in2<8> sl<60> vdd vss wl<8> / cell_PIM
XI25342 vss vss in1<16> in2<16> vss vdd vss wl<16> / cell_PIM
XI25341 vss vss in1<15> in2<15> vss vdd vss wl<15> / cell_PIM
XI25340 vss vss in1<17> in2<17> vss vdd vss wl<17> / cell_PIM
XI25339 vss vss in1<19> in2<19> vss vdd vss wl<19> / cell_PIM
XI25343 vss vss in1<13> in2<13> vss vdd vss wl<13> / cell_PIM
XI24688 bl<58> cbl<29> in1<9> in2<9> sl<58> vdd vss wl<9> / cell_PIM
XI25337 vss vss in1<21> in2<21> vss vdd vss wl<21> / cell_PIM
XI25336 vss vss in1<20> in2<20> vss vdd vss wl<20> / cell_PIM
XI25335 vss vss in1<24> in2<24> vss vdd vss wl<24> / cell_PIM
XI25334 vss vss in1<23> in2<23> vss vdd vss wl<23> / cell_PIM
XI25338 vss vss in1<18> in2<18> vss vdd vss wl<18> / cell_PIM
XI25332 vss vss in1<26> in2<26> vss vdd vss wl<26> / cell_PIM
XI25331 vss vss in1<25> in2<25> vss vdd vss wl<25> / cell_PIM
XI25330 vss vss in1<28> in2<28> vss vdd vss wl<28> / cell_PIM
XI25329 vss vss in1<27> in2<27> vss vdd vss wl<27> / cell_PIM
XI25333 vss vss in1<22> in2<22> vss vdd vss wl<22> / cell_PIM
XI25328 vss vss in1<31> in2<31> vss vdd vss wl<31> / cell_PIM
XI25327 vss vss in1<30> in2<30> vss vdd vss wl<30> / cell_PIM
XI25326 vss vss in1<29> in2<29> vss vdd vss wl<29> / cell_PIM
XI25325 vss vss in1<33> in2<33> vss vdd vss wl<33> / cell_PIM
XI25324 vss vss in1<32> in2<32> vss vdd vss wl<32> / cell_PIM
XI24678 bl<56> cbl<28> in1<9> in2<9> sl<56> vdd vss wl<9> / cell_PIM
XI25322 vss vss in1<34> in2<34> vss vdd vss wl<34> / cell_PIM
XI25321 vss vss in1<36> in2<36> vss vdd vss wl<36> / cell_PIM
XI25320 vss vss in1<38> in2<38> vss vdd vss wl<38> / cell_PIM
XI25319 vss vss in1<37> in2<37> vss vdd vss wl<37> / cell_PIM
XI25323 vss vss in1<35> in2<35> vss vdd vss wl<35> / cell_PIM
XI24668 bl<54> cbl<27> in1<9> in2<9> sl<54> vdd vss wl<9> / cell_PIM
XI25317 vss vss in1<39> in2<39> vss vdd vss wl<39> / cell_PIM
XI25316 vss vss in1<41> in2<41> vss vdd vss wl<41> / cell_PIM
XI25315 vss vss in1<43> in2<43> vss vdd vss wl<43> / cell_PIM
XI25314 vss vss in1<42> in2<42> vss vdd vss wl<42> / cell_PIM
XI25318 vss vss in1<40> in2<40> vss vdd vss wl<40> / cell_PIM
XI25312 vss vss in1<44> in2<44> vss vdd vss wl<44> / cell_PIM
XI25311 vss vss in1<47> in2<47> vss vdd vss wl<47> / cell_PIM
XI25310 vss vss in1<46> in2<46> vss vdd vss wl<46> / cell_PIM
XI25309 vss vss in1<50> in2<50> vss vdd vss wl<50> / cell_PIM
XI25313 vss vss in1<45> in2<45> vss vdd vss wl<45> / cell_PIM
XI25308 vss vss in1<49> in2<49> vss vdd vss wl<49> / cell_PIM
XI25307 vss vss in1<48> in2<48> vss vdd vss wl<48> / cell_PIM
XI25306 vss vss in1<52> in2<52> vss vdd vss wl<52> / cell_PIM
XI25305 vss vss in1<51> in2<51> vss vdd vss wl<51> / cell_PIM
XI25304 vss vss in1<55> in2<55> vss vdd vss wl<55> / cell_PIM
XI24658 bl<52> cbl<26> in1<8> in2<8> sl<52> vdd vss wl<8> / cell_PIM
XI25302 vss vss in1<53> in2<53> vss vdd vss wl<53> / cell_PIM
XI25301 vss vss in1<57> in2<57> vss vdd vss wl<57> / cell_PIM
XI25300 vss vss in1<56> in2<56> vss vdd vss wl<56> / cell_PIM
XI25299 vss vss in1<59> in2<59> vss vdd vss wl<59> / cell_PIM
XI25303 vss vss in1<54> in2<54> vss vdd vss wl<54> / cell_PIM
XI24648 bl<50> cbl<25> in1<9> in2<9> sl<50> vdd vss wl<9> / cell_PIM
XI25297 vss vss in1<60> in2<60> vss vdd vss wl<60> / cell_PIM
XI25296 vss vss in1<62> in2<62> vss vdd vss wl<62> / cell_PIM
XI25295 vss vss in1<61> in2<61> vss vdd vss wl<61> / cell_PIM
XI25294 vss vss in1<64> in2<64> vss vdd vss wl<64> / cell_PIM
XI25298 vss vss in1<58> in2<58> vss vdd vss wl<58> / cell_PIM
XI25292 vss vss in1<65> in2<65> vss vdd vss wl<65> / cell_PIM
XI25291 vss vss in1<67> in2<67> vss vdd vss wl<67> / cell_PIM
XI25290 vss vss in1<66> in2<66> vss vdd vss wl<66> / cell_PIM
XI25289 vss vss in1<69> in2<69> vss vdd vss wl<69> / cell_PIM
XI25293 vss vss in1<63> in2<63> vss vdd vss wl<63> / cell_PIM
XI25288 vss vss in1<68> in2<68> vss vdd vss wl<68> / cell_PIM
XI25287 vss vss in1<70> in2<70> vss vdd vss wl<70> / cell_PIM
XI25286 vss vss in1<71> in2<71> vss vdd vss wl<71> / cell_PIM
XI25285 vss vss in1<74> in2<74> vss vdd vss wl<74> / cell_PIM
XI25284 vss vss in1<73> in2<73> vss vdd vss wl<73> / cell_PIM
XI24638 bl<48> cbl<24> in1<8> in2<8> sl<48> vdd vss wl<8> / cell_PIM
XI25282 vss vss in1<75> in2<75> vss vdd vss wl<75> / cell_PIM
XI25281 vss vss in1<76> in2<76> vss vdd vss wl<76> / cell_PIM
XI25280 vss vss in1<79> in2<79> vss vdd vss wl<79> / cell_PIM
XI25279 vss vss in1<78> in2<78> vss vdd vss wl<78> / cell_PIM
XI25283 vss vss in1<72> in2<72> vss vdd vss wl<72> / cell_PIM
XI24628 bl<46> cbl<23> in1<9> in2<9> sl<46> vdd vss wl<9> / cell_PIM
XI25277 vss vss in1<80> in2<80> vss vdd vss wl<80> / cell_PIM
XI25276 vss vss in1<81> in2<81> vss vdd vss wl<81> / cell_PIM
XI25275 vss vss in1<83> in2<83> vss vdd vss wl<83> / cell_PIM
XI25274 vss vss in1<82> in2<82> vss vdd vss wl<82> / cell_PIM
XI25278 vss vss in1<77> in2<77> vss vdd vss wl<77> / cell_PIM
XI25272 vss vss in1<86> in2<86> vss vdd vss wl<86> / cell_PIM
XI25271 vss vss in1<85> in2<85> vss vdd vss wl<85> / cell_PIM
XI25270 vss vss in1<88> in2<88> vss vdd vss wl<88> / cell_PIM
XI25269 vss vss in1<87> in2<87> vss vdd vss wl<87> / cell_PIM
XI25273 vss vss in1<84> in2<84> vss vdd vss wl<84> / cell_PIM
XI25268 vss vss in1<89> in2<89> vss vdd vss wl<89> / cell_PIM
XI25267 vss vss in1<91> in2<91> vss vdd vss wl<91> / cell_PIM
XI25266 vss vss in1<90> in2<90> vss vdd vss wl<90> / cell_PIM
XI25265 vss vss in1<93> in2<93> vss vdd vss wl<93> / cell_PIM
XI25264 vss vss in1<92> in2<92> vss vdd vss wl<92> / cell_PIM
XI24618 bl<44> cbl<22> in1<8> in2<8> sl<44> vdd vss wl<8> / cell_PIM
XI25262 vss vss in1<95> in2<95> vss vdd vss wl<95> / cell_PIM
XI25261 vss vss in1<98> in2<98> vss vdd vss wl<98> / cell_PIM
XI25260 vss vss in1<97> in2<97> vss vdd vss wl<97> / cell_PIM
XI25259 vss vss in1<96> in2<96> vss vdd vss wl<96> / cell_PIM
XI25263 vss vss in1<94> in2<94> vss vdd vss wl<94> / cell_PIM
XI24608 bl<42> cbl<21> in1<9> in2<9> sl<42> vdd vss wl<9> / cell_PIM
XI25257 vss vss in1<100> in2<100> vss vdd vss wl<100> / cell_PIM
XI25256 vss vss in1<103> in2<103> vss vdd vss wl<103> / cell_PIM
XI25255 vss vss in1<102> in2<102> vss vdd vss wl<102> / cell_PIM
XI25254 vss vss in1<101> in2<101> vss vdd vss wl<101> / cell_PIM
XI25258 vss vss in1<99> in2<99> vss vdd vss wl<99> / cell_PIM
XI25252 vss vss in1<105> in2<105> vss vdd vss wl<105> / cell_PIM
XI25251 vss vss in1<107> in2<107> vss vdd vss wl<107> / cell_PIM
XI25250 vss vss in1<106> in2<106> vss vdd vss wl<106> / cell_PIM
XI25249 vss vss in1<108> in2<108> vss vdd vss wl<108> / cell_PIM
XI25253 vss vss in1<104> in2<104> vss vdd vss wl<104> / cell_PIM
XI25248 vss vss in1<109> in2<109> vss vdd vss wl<109> / cell_PIM
XI25247 vss vss in1<110> in2<110> vss vdd vss wl<110> / cell_PIM
XI25246 vss vss in1<112> in2<112> vss vdd vss wl<112> / cell_PIM
XI25245 vss vss in1<111> in2<111> vss vdd vss wl<111> / cell_PIM
XI25244 vss vss in1<113> in2<113> vss vdd vss wl<113> / cell_PIM
XI24598 bl<40> cbl<20> in1<9> in2<9> sl<40> vdd vss wl<9> / cell_PIM
XI25242 vss vss in1<115> in2<115> vss vdd vss wl<115> / cell_PIM
XI25241 vss vss in1<117> in2<117> vss vdd vss wl<117> / cell_PIM
XI25240 vss vss in1<116> in2<116> vss vdd vss wl<116> / cell_PIM
XI25239 vss vss in1<118> in2<118> vss vdd vss wl<118> / cell_PIM
XI25243 vss vss in1<114> in2<114> vss vdd vss wl<114> / cell_PIM
XI24588 bl<38> cbl<19> in1<9> in2<9> sl<38> vdd vss wl<9> / cell_PIM
XI25237 vss vss in1<122> in2<122> vss vdd vss wl<122> / cell_PIM
XI25236 vss vss in1<121> in2<121> vss vdd vss wl<121> / cell_PIM
XI25235 vss vss in1<120> in2<120> vss vdd vss wl<120> / cell_PIM
XI25234 vss vss in1<123> in2<123> vss vdd vss wl<123> / cell_PIM
XI25238 vss vss in1<119> in2<119> vss vdd vss wl<119> / cell_PIM
XI25232 vss vss in1<127> in2<127> vss vdd vss wl<127> / cell_PIM
XI25231 vss vss in1<126> in2<126> vss vdd vss wl<126> / cell_PIM
XI25230 vss vss in1<125> in2<125> vss vdd vss wl<125> / cell_PIM
XI25229 vss vss in1<124> in2<124> vss vdd vss wl<124> / cell_PIM
XI25233 vss vss vdd vdd vss vdd vss vss / cell_PIM
XI24578 bl<36> cbl<18> in1<8> in2<8> sl<36> vdd vss wl<8> / cell_PIM
XI24568 bl<34> cbl<17> in1<9> in2<9> sl<34> vdd vss wl<9> / cell_PIM
XI24558 bl<32> cbl<16> in1<8> in2<8> sl<32> vdd vss wl<8> / cell_PIM
XI24548 bl<62> cbl<31> in1<14> in2<14> sl<62> vdd vss wl<14> / cell_PIM
XI24538 bl<60> cbl<30> in1<13> in2<13> sl<60> vdd vss wl<13> / cell_PIM
XI24528 bl<58> cbl<29> in1<14> in2<14> sl<58> vdd vss wl<14> / cell_PIM
XI24518 bl<56> cbl<28> in1<14> in2<14> sl<56> vdd vss wl<14> / cell_PIM
XI24508 bl<54> cbl<27> in1<14> in2<14> sl<54> vdd vss wl<14> / cell_PIM
XI24498 bl<52> cbl<26> in1<13> in2<13> sl<52> vdd vss wl<13> / cell_PIM
XI24488 bl<50> cbl<25> in1<14> in2<14> sl<50> vdd vss wl<14> / cell_PIM
XI24478 bl<48> cbl<24> in1<13> in2<13> sl<48> vdd vss wl<13> / cell_PIM
XI24468 bl<46> cbl<23> in1<14> in2<14> sl<46> vdd vss wl<14> / cell_PIM
XI24458 bl<44> cbl<22> in1<13> in2<13> sl<44> vdd vss wl<13> / cell_PIM
XI24448 bl<42> cbl<21> in1<14> in2<14> sl<42> vdd vss wl<14> / cell_PIM
XI25097 bl<62> cbl<31> vdd vdd sl<62> vdd vss vss / cell_PIM
XI25095 bl<60> cbl<30> vdd vdd sl<60> vdd vss vss / cell_PIM
XI25091 bl<56> cbl<28> vdd vdd sl<56> vdd vss vss / cell_PIM
XI25089 bl<54> cbl<27> vdd vdd sl<54> vdd vss vss / cell_PIM
XI25093 bl<58> cbl<29> vdd vdd sl<58> vdd vss vss / cell_PIM
XI25087 bl<52> cbl<26> vdd vdd sl<52> vdd vss vss / cell_PIM
XI25085 bl<50> cbl<25> vdd vdd sl<50> vdd vss vss / cell_PIM
XI24438 bl<40> cbl<20> in1<14> in2<14> sl<40> vdd vss wl<14> / cell_PIM
XI25081 bl<46> cbl<23> vdd vdd sl<46> vdd vss vss / cell_PIM
XI25079 bl<44> cbl<22> vdd vdd sl<44> vdd vss vss / cell_PIM
XI25083 bl<48> cbl<24> vdd vdd sl<48> vdd vss vss / cell_PIM
XI24428 bl<38> cbl<19> in1<14> in2<14> sl<38> vdd vss wl<14> / cell_PIM
XI25077 bl<42> cbl<21> vdd vdd sl<42> vdd vss vss / cell_PIM
XI25075 bl<40> cbl<20> vdd vdd sl<40> vdd vss vss / cell_PIM
XI25071 bl<36> cbl<18> vdd vdd sl<36> vdd vss vss / cell_PIM
XI25069 bl<34> cbl<17> vdd vdd sl<34> vdd vss vss / cell_PIM
XI25073 bl<38> cbl<19> vdd vdd sl<38> vdd vss vss / cell_PIM
XI25067 bl<32> cbl<16> vdd vdd sl<32> vdd vss vss / cell_PIM
XI25065 bl<30> cbl<15> vdd vdd sl<30> vdd vss vss / cell_PIM
XI24418 bl<36> cbl<18> in1<13> in2<13> sl<36> vdd vss wl<13> / cell_PIM
XI25061 bl<26> cbl<13> vdd vdd sl<26> vdd vss vss / cell_PIM
XI25059 bl<24> cbl<12> vdd vdd sl<24> vdd vss vss / cell_PIM
XI25063 bl<28> cbl<14> vdd vdd sl<28> vdd vss vss / cell_PIM
XI24408 bl<34> cbl<17> in1<14> in2<14> sl<34> vdd vss wl<14> / cell_PIM
XI25057 bl<22> cbl<11> vdd vdd sl<22> vdd vss vss / cell_PIM
XI25055 bl<20> cbl<10> vdd vdd sl<20> vdd vss vss / cell_PIM
XI25051 bl<16> cbl<8> vdd vdd sl<16> vdd vss vss / cell_PIM
XI25049 bl<14> cbl<7> vdd vdd sl<14> vdd vss vss / cell_PIM
XI25053 bl<18> cbl<9> vdd vdd sl<18> vdd vss vss / cell_PIM
XI25047 bl<12> cbl<6> vdd vdd sl<12> vdd vss vss / cell_PIM
XI25045 bl<10> cbl<5> vdd vdd sl<10> vdd vss vss / cell_PIM
XI24398 bl<32> cbl<16> in1<13> in2<13> sl<32> vdd vss wl<13> / cell_PIM
XI25041 bl<6> cbl<3> vdd vdd sl<6> vdd vss vss / cell_PIM
XI25039 bl<4> cbl<2> vdd vdd sl<4> vdd vss vss / cell_PIM
XI25043 bl<8> cbl<4> vdd vdd sl<8> vdd vss vss / cell_PIM
XI24388 bl<62> cbl<31> in1<21> in2<21> sl<62> vdd vss wl<21> / cell_PIM
XI25037 bl<2> cbl<1> vdd vdd sl<2> vdd vss vss / cell_PIM
XI25035 bl<0> cbl<0> vdd vdd sl<0> vdd vss vss / cell_PIM
XI22883 bl<62> cbl<31> in1<67> in2<67> sl<62> vdd vss wl<67> / cell_PIM
XI23403 bl<44> cbl<22> in1<47> in2<47> sl<44> vdd vss wl<47> / cell_PIM
XI23402 bl<44> cbl<22> in1<46> in2<46> sl<44> vdd vss wl<46> / cell_PIM
XI23401 bl<44> cbl<22> in1<50> in2<50> sl<44> vdd vss wl<50> / cell_PIM
XI24051 bl<52> cbl<26> in1<28> in2<28> sl<52> vdd vss wl<28> / cell_PIM
XI24050 bl<52> cbl<26> in1<27> in2<27> sl<52> vdd vss wl<27> / cell_PIM
XI24049 bl<52> cbl<26> in1<31> in2<31> sl<52> vdd vss wl<31> / cell_PIM
XI24699 bl<60> cbl<30> in1<9> in2<9> sl<60> vdd vss wl<9> / cell_PIM
XI24697 bl<60> cbl<30> in1<12> in2<12> sl<60> vdd vss wl<12> / cell_PIM
XI24696 bl<60> cbl<30> in1<11> in2<11> sl<60> vdd vss wl<11> / cell_PIM
XI24695 bl<60> cbl<30> in1<10> in2<10> sl<60> vdd vss wl<10> / cell_PIM
XI24048 bl<52> cbl<26> in1<30> in2<30> sl<52> vdd vss wl<30> / cell_PIM
XI24047 bl<52> cbl<26> in1<29> in2<29> sl<52> vdd vss wl<29> / cell_PIM
XI23400 bl<44> cbl<22> in1<49> in2<49> sl<44> vdd vss wl<49> / cell_PIM
XI23399 bl<44> cbl<22> in1<48> in2<48> sl<44> vdd vss wl<48> / cell_PIM
XI22873 bl<60> cbl<30> in1<65> in2<65> sl<60> vdd vss wl<65> / cell_PIM
XI23393 bl<42> cbl<21> in1<46> in2<46> sl<42> vdd vss wl<46> / cell_PIM
XI24041 bl<50> cbl<25> in1<27> in2<27> sl<50> vdd vss wl<27> / cell_PIM
XI24040 bl<50> cbl<25> in1<28> in2<28> sl<50> vdd vss wl<28> / cell_PIM
XI24039 bl<50> cbl<25> in1<30> in2<30> sl<50> vdd vss wl<30> / cell_PIM
XI24689 bl<58> cbl<29> in1<8> in2<8> sl<58> vdd vss wl<8> / cell_PIM
XI23392 bl<42> cbl<21> in1<47> in2<47> sl<42> vdd vss wl<47> / cell_PIM
XI23391 bl<42> cbl<21> in1<49> in2<49> sl<42> vdd vss wl<49> / cell_PIM
XI23390 bl<42> cbl<21> in1<50> in2<50> sl<42> vdd vss wl<50> / cell_PIM
XI23389 bl<42> cbl<21> in1<48> in2<48> sl<42> vdd vss wl<48> / cell_PIM
XI24038 bl<50> cbl<25> in1<31> in2<31> sl<50> vdd vss wl<31> / cell_PIM
XI24037 bl<50> cbl<25> in1<29> in2<29> sl<50> vdd vss wl<29> / cell_PIM
XI24687 bl<58> cbl<29> in1<11> in2<11> sl<58> vdd vss wl<11> / cell_PIM
XI24686 bl<58> cbl<29> in1<12> in2<12> sl<58> vdd vss wl<12> / cell_PIM
XI24685 bl<58> cbl<29> in1<10> in2<10> sl<58> vdd vss wl<10> / cell_PIM
XI22863 bl<58> cbl<29> in1<67> in2<67> sl<58> vdd vss wl<67> / cell_PIM
XI24031 bl<48> cbl<24> in1<28> in2<28> sl<48> vdd vss wl<28> / cell_PIM
XI24030 bl<48> cbl<24> in1<27> in2<27> sl<48> vdd vss wl<27> / cell_PIM
XI24029 bl<48> cbl<24> in1<31> in2<31> sl<48> vdd vss wl<31> / cell_PIM
XI24679 bl<56> cbl<28> in1<8> in2<8> sl<56> vdd vss wl<8> / cell_PIM
XI24677 bl<56> cbl<28> in1<11> in2<11> sl<56> vdd vss wl<11> / cell_PIM
XI24676 bl<56> cbl<28> in1<12> in2<12> sl<56> vdd vss wl<12> / cell_PIM
XI24675 bl<56> cbl<28> in1<10> in2<10> sl<56> vdd vss wl<10> / cell_PIM
XI24028 bl<48> cbl<24> in1<30> in2<30> sl<48> vdd vss wl<30> / cell_PIM
XI24027 bl<48> cbl<24> in1<29> in2<29> sl<48> vdd vss wl<29> / cell_PIM
XI23383 bl<40> cbl<20> in1<46> in2<46> sl<40> vdd vss wl<46> / cell_PIM
XI23382 bl<40> cbl<20> in1<47> in2<47> sl<40> vdd vss wl<47> / cell_PIM
XI23381 bl<40> cbl<20> in1<49> in2<49> sl<40> vdd vss wl<49> / cell_PIM
XI22853 bl<56> cbl<28> in1<67> in2<67> sl<56> vdd vss wl<67> / cell_PIM
XI23380 bl<40> cbl<20> in1<50> in2<50> sl<40> vdd vss wl<50> / cell_PIM
XI23379 bl<40> cbl<20> in1<48> in2<48> sl<40> vdd vss wl<48> / cell_PIM
XI24021 bl<46> cbl<23> in1<27> in2<27> sl<46> vdd vss wl<27> / cell_PIM
XI24020 bl<46> cbl<23> in1<28> in2<28> sl<46> vdd vss wl<28> / cell_PIM
XI24019 bl<46> cbl<23> in1<30> in2<30> sl<46> vdd vss wl<30> / cell_PIM
XI24669 bl<54> cbl<27> in1<8> in2<8> sl<54> vdd vss wl<8> / cell_PIM
XI23373 bl<38> cbl<19> in1<46> in2<46> sl<38> vdd vss wl<46> / cell_PIM
XI24018 bl<46> cbl<23> in1<31> in2<31> sl<46> vdd vss wl<31> / cell_PIM
XI24017 bl<46> cbl<23> in1<29> in2<29> sl<46> vdd vss wl<29> / cell_PIM
XI24667 bl<54> cbl<27> in1<11> in2<11> sl<54> vdd vss wl<11> / cell_PIM
XI24666 bl<54> cbl<27> in1<12> in2<12> sl<54> vdd vss wl<12> / cell_PIM
XI24665 bl<54> cbl<27> in1<10> in2<10> sl<54> vdd vss wl<10> / cell_PIM
XI22843 bl<54> cbl<27> in1<67> in2<67> sl<54> vdd vss wl<67> / cell_PIM
XI23372 bl<38> cbl<19> in1<47> in2<47> sl<38> vdd vss wl<47> / cell_PIM
XI23371 bl<38> cbl<19> in1<49> in2<49> sl<38> vdd vss wl<49> / cell_PIM
XI23370 bl<38> cbl<19> in1<50> in2<50> sl<38> vdd vss wl<50> / cell_PIM
XI23369 bl<38> cbl<19> in1<48> in2<48> sl<38> vdd vss wl<48> / cell_PIM
XI24011 bl<44> cbl<22> in1<28> in2<28> sl<44> vdd vss wl<28> / cell_PIM
XI24010 bl<44> cbl<22> in1<27> in2<27> sl<44> vdd vss wl<27> / cell_PIM
XI24009 bl<44> cbl<22> in1<31> in2<31> sl<44> vdd vss wl<31> / cell_PIM
XI24659 bl<52> cbl<26> in1<9> in2<9> sl<52> vdd vss wl<9> / cell_PIM
XI24657 bl<52> cbl<26> in1<12> in2<12> sl<52> vdd vss wl<12> / cell_PIM
XI24656 bl<52> cbl<26> in1<11> in2<11> sl<52> vdd vss wl<11> / cell_PIM
XI24655 bl<52> cbl<26> in1<10> in2<10> sl<52> vdd vss wl<10> / cell_PIM
XI24008 bl<44> cbl<22> in1<30> in2<30> sl<44> vdd vss wl<30> / cell_PIM
XI24007 bl<44> cbl<22> in1<29> in2<29> sl<44> vdd vss wl<29> / cell_PIM
XI22833 bl<52> cbl<26> in1<65> in2<65> sl<52> vdd vss wl<65> / cell_PIM
XI23363 bl<36> cbl<18> in1<47> in2<47> sl<36> vdd vss wl<47> / cell_PIM
XI23362 bl<36> cbl<18> in1<46> in2<46> sl<36> vdd vss wl<46> / cell_PIM
XI23361 bl<36> cbl<18> in1<50> in2<50> sl<36> vdd vss wl<50> / cell_PIM
XI24001 bl<42> cbl<21> in1<27> in2<27> sl<42> vdd vss wl<27> / cell_PIM
XI24000 bl<42> cbl<21> in1<28> in2<28> sl<42> vdd vss wl<28> / cell_PIM
XI23999 bl<42> cbl<21> in1<30> in2<30> sl<42> vdd vss wl<30> / cell_PIM
XI24649 bl<50> cbl<25> in1<8> in2<8> sl<50> vdd vss wl<8> / cell_PIM
XI23360 bl<36> cbl<18> in1<49> in2<49> sl<36> vdd vss wl<49> / cell_PIM
XI23359 bl<36> cbl<18> in1<48> in2<48> sl<36> vdd vss wl<48> / cell_PIM
XI23998 bl<42> cbl<21> in1<31> in2<31> sl<42> vdd vss wl<31> / cell_PIM
XI23997 bl<42> cbl<21> in1<29> in2<29> sl<42> vdd vss wl<29> / cell_PIM
XI24647 bl<50> cbl<25> in1<11> in2<11> sl<50> vdd vss wl<11> / cell_PIM
XI24646 bl<50> cbl<25> in1<12> in2<12> sl<50> vdd vss wl<12> / cell_PIM
XI24645 bl<50> cbl<25> in1<10> in2<10> sl<50> vdd vss wl<10> / cell_PIM
XI22823 bl<50> cbl<25> in1<67> in2<67> sl<50> vdd vss wl<67> / cell_PIM
XI23353 bl<34> cbl<17> in1<46> in2<46> sl<34> vdd vss wl<46> / cell_PIM
XI23991 bl<40> cbl<20> in1<27> in2<27> sl<40> vdd vss wl<27> / cell_PIM
XI23990 bl<40> cbl<20> in1<28> in2<28> sl<40> vdd vss wl<28> / cell_PIM
XI23989 bl<40> cbl<20> in1<30> in2<30> sl<40> vdd vss wl<30> / cell_PIM
XI24639 bl<48> cbl<24> in1<9> in2<9> sl<48> vdd vss wl<9> / cell_PIM
XI24637 bl<48> cbl<24> in1<12> in2<12> sl<48> vdd vss wl<12> / cell_PIM
XI24636 bl<48> cbl<24> in1<11> in2<11> sl<48> vdd vss wl<11> / cell_PIM
XI24635 bl<48> cbl<24> in1<10> in2<10> sl<48> vdd vss wl<10> / cell_PIM
XI23988 bl<40> cbl<20> in1<31> in2<31> sl<40> vdd vss wl<31> / cell_PIM
XI23987 bl<40> cbl<20> in1<29> in2<29> sl<40> vdd vss wl<29> / cell_PIM
XI23352 bl<34> cbl<17> in1<47> in2<47> sl<34> vdd vss wl<47> / cell_PIM
XI23351 bl<34> cbl<17> in1<49> in2<49> sl<34> vdd vss wl<49> / cell_PIM
XI23350 bl<34> cbl<17> in1<50> in2<50> sl<34> vdd vss wl<50> / cell_PIM
XI23349 bl<34> cbl<17> in1<48> in2<48> sl<34> vdd vss wl<48> / cell_PIM
XI22813 bl<48> cbl<24> in1<65> in2<65> sl<48> vdd vss wl<65> / cell_PIM
XI23981 bl<38> cbl<19> in1<27> in2<27> sl<38> vdd vss wl<27> / cell_PIM
XI23980 bl<38> cbl<19> in1<28> in2<28> sl<38> vdd vss wl<28> / cell_PIM
XI23979 bl<38> cbl<19> in1<30> in2<30> sl<38> vdd vss wl<30> / cell_PIM
XI24629 bl<46> cbl<23> in1<8> in2<8> sl<46> vdd vss wl<8> / cell_PIM
XI23343 bl<32> cbl<16> in1<47> in2<47> sl<32> vdd vss wl<47> / cell_PIM
XI23342 bl<32> cbl<16> in1<46> in2<46> sl<32> vdd vss wl<46> / cell_PIM
XI23341 bl<32> cbl<16> in1<50> in2<50> sl<32> vdd vss wl<50> / cell_PIM
XI23978 bl<38> cbl<19> in1<31> in2<31> sl<38> vdd vss wl<31> / cell_PIM
XI23977 bl<38> cbl<19> in1<29> in2<29> sl<38> vdd vss wl<29> / cell_PIM
XI24627 bl<46> cbl<23> in1<11> in2<11> sl<46> vdd vss wl<11> / cell_PIM
XI24626 bl<46> cbl<23> in1<12> in2<12> sl<46> vdd vss wl<12> / cell_PIM
XI24625 bl<46> cbl<23> in1<10> in2<10> sl<46> vdd vss wl<10> / cell_PIM
XI22803 bl<46> cbl<23> in1<67> in2<67> sl<46> vdd vss wl<67> / cell_PIM
XI23340 bl<32> cbl<16> in1<49> in2<49> sl<32> vdd vss wl<49> / cell_PIM
XI23339 bl<32> cbl<16> in1<48> in2<48> sl<32> vdd vss wl<48> / cell_PIM
XI23971 bl<36> cbl<18> in1<28> in2<28> sl<36> vdd vss wl<28> / cell_PIM
XI23970 bl<36> cbl<18> in1<27> in2<27> sl<36> vdd vss wl<27> / cell_PIM
XI23969 bl<36> cbl<18> in1<31> in2<31> sl<36> vdd vss wl<31> / cell_PIM
XI24619 bl<44> cbl<22> in1<9> in2<9> sl<44> vdd vss wl<9> / cell_PIM
XI24617 bl<44> cbl<22> in1<12> in2<12> sl<44> vdd vss wl<12> / cell_PIM
XI24616 bl<44> cbl<22> in1<11> in2<11> sl<44> vdd vss wl<11> / cell_PIM
XI24615 bl<44> cbl<22> in1<10> in2<10> sl<44> vdd vss wl<10> / cell_PIM
XI23968 bl<36> cbl<18> in1<30> in2<30> sl<36> vdd vss wl<30> / cell_PIM
XI23967 bl<36> cbl<18> in1<29> in2<29> sl<36> vdd vss wl<29> / cell_PIM
XI23333 bl<62> cbl<31> in1<51> in2<51> sl<62> vdd vss wl<51> / cell_PIM
XI22793 bl<44> cbl<22> in1<65> in2<65> sl<44> vdd vss wl<65> / cell_PIM
XI23332 bl<62> cbl<31> in1<52> in2<52> sl<62> vdd vss wl<52> / cell_PIM
XI23331 bl<62> cbl<31> in1<54> in2<54> sl<62> vdd vss wl<54> / cell_PIM
XI23330 bl<62> cbl<31> in1<55> in2<55> sl<62> vdd vss wl<55> / cell_PIM
XI23329 bl<62> cbl<31> in1<53> in2<53> sl<62> vdd vss wl<53> / cell_PIM
XI23961 bl<34> cbl<17> in1<27> in2<27> sl<34> vdd vss wl<27> / cell_PIM
XI23960 bl<34> cbl<17> in1<28> in2<28> sl<34> vdd vss wl<28> / cell_PIM
XI23959 bl<34> cbl<17> in1<30> in2<30> sl<34> vdd vss wl<30> / cell_PIM
XI24609 bl<42> cbl<21> in1<8> in2<8> sl<42> vdd vss wl<8> / cell_PIM
XI23958 bl<34> cbl<17> in1<31> in2<31> sl<34> vdd vss wl<31> / cell_PIM
XI23957 bl<34> cbl<17> in1<29> in2<29> sl<34> vdd vss wl<29> / cell_PIM
XI24607 bl<42> cbl<21> in1<11> in2<11> sl<42> vdd vss wl<11> / cell_PIM
XI24606 bl<42> cbl<21> in1<12> in2<12> sl<42> vdd vss wl<12> / cell_PIM
XI24605 bl<42> cbl<21> in1<10> in2<10> sl<42> vdd vss wl<10> / cell_PIM
XI22783 bl<42> cbl<21> in1<67> in2<67> sl<42> vdd vss wl<67> / cell_PIM
XI23323 bl<60> cbl<30> in1<52> in2<52> sl<60> vdd vss wl<52> / cell_PIM
XI23322 bl<60> cbl<30> in1<51> in2<51> sl<60> vdd vss wl<51> / cell_PIM
XI23321 bl<60> cbl<30> in1<55> in2<55> sl<60> vdd vss wl<55> / cell_PIM
XI23951 bl<32> cbl<16> in1<28> in2<28> sl<32> vdd vss wl<28> / cell_PIM
XI23950 bl<32> cbl<16> in1<27> in2<27> sl<32> vdd vss wl<27> / cell_PIM
XI23949 bl<32> cbl<16> in1<31> in2<31> sl<32> vdd vss wl<31> / cell_PIM
XI24599 bl<40> cbl<20> in1<8> in2<8> sl<40> vdd vss wl<8> / cell_PIM
XI24597 bl<40> cbl<20> in1<11> in2<11> sl<40> vdd vss wl<11> / cell_PIM
XI24596 bl<40> cbl<20> in1<12> in2<12> sl<40> vdd vss wl<12> / cell_PIM
XI24595 bl<40> cbl<20> in1<10> in2<10> sl<40> vdd vss wl<10> / cell_PIM
XI23948 bl<32> cbl<16> in1<30> in2<30> sl<32> vdd vss wl<30> / cell_PIM
XI23947 bl<32> cbl<16> in1<29> in2<29> sl<32> vdd vss wl<29> / cell_PIM
XI23320 bl<60> cbl<30> in1<54> in2<54> sl<60> vdd vss wl<54> / cell_PIM
XI23319 bl<60> cbl<30> in1<53> in2<53> sl<60> vdd vss wl<53> / cell_PIM
XI22773 bl<40> cbl<20> in1<67> in2<67> sl<40> vdd vss wl<67> / cell_PIM
XI23313 bl<58> cbl<29> in1<51> in2<51> sl<58> vdd vss wl<51> / cell_PIM
XI23941 bl<62> cbl<31> in1<32> in2<32> sl<62> vdd vss wl<32> / cell_PIM
XI23940 bl<62> cbl<31> in1<33> in2<33> sl<62> vdd vss wl<33> / cell_PIM
XI23939 bl<62> cbl<31> in1<35> in2<35> sl<62> vdd vss wl<35> / cell_PIM
XI24589 bl<38> cbl<19> in1<8> in2<8> sl<38> vdd vss wl<8> / cell_PIM
XI23312 bl<58> cbl<29> in1<52> in2<52> sl<58> vdd vss wl<52> / cell_PIM
XI23311 bl<58> cbl<29> in1<54> in2<54> sl<58> vdd vss wl<54> / cell_PIM
XI23310 bl<58> cbl<29> in1<55> in2<55> sl<58> vdd vss wl<55> / cell_PIM
XI23309 bl<58> cbl<29> in1<53> in2<53> sl<58> vdd vss wl<53> / cell_PIM
XI23938 bl<62> cbl<31> in1<36> in2<36> sl<62> vdd vss wl<36> / cell_PIM
XI23937 bl<62> cbl<31> in1<34> in2<34> sl<62> vdd vss wl<34> / cell_PIM
XI24587 bl<38> cbl<19> in1<11> in2<11> sl<38> vdd vss wl<11> / cell_PIM
XI24586 bl<38> cbl<19> in1<12> in2<12> sl<38> vdd vss wl<12> / cell_PIM
XI24585 bl<38> cbl<19> in1<10> in2<10> sl<38> vdd vss wl<10> / cell_PIM
XI22763 bl<38> cbl<19> in1<67> in2<67> sl<38> vdd vss wl<67> / cell_PIM
XI23931 bl<60> cbl<30> in1<33> in2<33> sl<60> vdd vss wl<33> / cell_PIM
XI23930 bl<60> cbl<30> in1<32> in2<32> sl<60> vdd vss wl<32> / cell_PIM
XI23929 bl<60> cbl<30> in1<36> in2<36> sl<60> vdd vss wl<36> / cell_PIM
XI24579 bl<36> cbl<18> in1<9> in2<9> sl<36> vdd vss wl<9> / cell_PIM
XI24577 bl<36> cbl<18> in1<12> in2<12> sl<36> vdd vss wl<12> / cell_PIM
XI24576 bl<36> cbl<18> in1<11> in2<11> sl<36> vdd vss wl<11> / cell_PIM
XI24575 bl<36> cbl<18> in1<10> in2<10> sl<36> vdd vss wl<10> / cell_PIM
XI23928 bl<60> cbl<30> in1<35> in2<35> sl<60> vdd vss wl<35> / cell_PIM
XI23927 bl<60> cbl<30> in1<34> in2<34> sl<60> vdd vss wl<34> / cell_PIM
XI23303 bl<56> cbl<28> in1<51> in2<51> sl<56> vdd vss wl<51> / cell_PIM
XI23302 bl<56> cbl<28> in1<52> in2<52> sl<56> vdd vss wl<52> / cell_PIM
XI23301 bl<56> cbl<28> in1<54> in2<54> sl<56> vdd vss wl<54> / cell_PIM
XI22753 bl<36> cbl<18> in1<65> in2<65> sl<36> vdd vss wl<65> / cell_PIM
XI23300 bl<56> cbl<28> in1<55> in2<55> sl<56> vdd vss wl<55> / cell_PIM
XI23299 bl<56> cbl<28> in1<53> in2<53> sl<56> vdd vss wl<53> / cell_PIM
XI23921 bl<58> cbl<29> in1<32> in2<32> sl<58> vdd vss wl<32> / cell_PIM
XI23920 bl<58> cbl<29> in1<33> in2<33> sl<58> vdd vss wl<33> / cell_PIM
XI23919 bl<58> cbl<29> in1<35> in2<35> sl<58> vdd vss wl<35> / cell_PIM
XI24569 bl<34> cbl<17> in1<8> in2<8> sl<34> vdd vss wl<8> / cell_PIM
XI23293 bl<54> cbl<27> in1<51> in2<51> sl<54> vdd vss wl<51> / cell_PIM
XI23918 bl<58> cbl<29> in1<36> in2<36> sl<58> vdd vss wl<36> / cell_PIM
XI23917 bl<58> cbl<29> in1<34> in2<34> sl<58> vdd vss wl<34> / cell_PIM
XI24567 bl<34> cbl<17> in1<11> in2<11> sl<34> vdd vss wl<11> / cell_PIM
XI24566 bl<34> cbl<17> in1<12> in2<12> sl<34> vdd vss wl<12> / cell_PIM
XI24565 bl<34> cbl<17> in1<10> in2<10> sl<34> vdd vss wl<10> / cell_PIM
XI22743 bl<34> cbl<17> in1<67> in2<67> sl<34> vdd vss wl<67> / cell_PIM
XI23292 bl<54> cbl<27> in1<52> in2<52> sl<54> vdd vss wl<52> / cell_PIM
XI23291 bl<54> cbl<27> in1<54> in2<54> sl<54> vdd vss wl<54> / cell_PIM
XI23290 bl<54> cbl<27> in1<55> in2<55> sl<54> vdd vss wl<55> / cell_PIM
XI23289 bl<54> cbl<27> in1<53> in2<53> sl<54> vdd vss wl<53> / cell_PIM
XI23911 bl<56> cbl<28> in1<32> in2<32> sl<56> vdd vss wl<32> / cell_PIM
XI23910 bl<56> cbl<28> in1<33> in2<33> sl<56> vdd vss wl<33> / cell_PIM
XI23909 bl<56> cbl<28> in1<35> in2<35> sl<56> vdd vss wl<35> / cell_PIM
XI24559 bl<32> cbl<16> in1<9> in2<9> sl<32> vdd vss wl<9> / cell_PIM
XI24557 bl<32> cbl<16> in1<12> in2<12> sl<32> vdd vss wl<12> / cell_PIM
XI24556 bl<32> cbl<16> in1<11> in2<11> sl<32> vdd vss wl<11> / cell_PIM
XI24555 bl<32> cbl<16> in1<10> in2<10> sl<32> vdd vss wl<10> / cell_PIM
XI23908 bl<56> cbl<28> in1<36> in2<36> sl<56> vdd vss wl<36> / cell_PIM
XI23907 bl<56> cbl<28> in1<34> in2<34> sl<56> vdd vss wl<34> / cell_PIM
XI22733 bl<32> cbl<16> in1<65> in2<65> sl<32> vdd vss wl<65> / cell_PIM
XI23283 bl<52> cbl<26> in1<52> in2<52> sl<52> vdd vss wl<52> / cell_PIM
XI23282 bl<52> cbl<26> in1<51> in2<51> sl<52> vdd vss wl<51> / cell_PIM
XI23281 bl<52> cbl<26> in1<55> in2<55> sl<52> vdd vss wl<55> / cell_PIM
XI23901 bl<54> cbl<27> in1<32> in2<32> sl<54> vdd vss wl<32> / cell_PIM
XI23900 bl<54> cbl<27> in1<33> in2<33> sl<54> vdd vss wl<33> / cell_PIM
XI23899 bl<54> cbl<27> in1<35> in2<35> sl<54> vdd vss wl<35> / cell_PIM
XI24549 bl<62> cbl<31> in1<13> in2<13> sl<62> vdd vss wl<13> / cell_PIM
XI23280 bl<52> cbl<26> in1<54> in2<54> sl<52> vdd vss wl<54> / cell_PIM
XI23279 bl<52> cbl<26> in1<53> in2<53> sl<52> vdd vss wl<53> / cell_PIM
XI23898 bl<54> cbl<27> in1<36> in2<36> sl<54> vdd vss wl<36> / cell_PIM
XI23897 bl<54> cbl<27> in1<34> in2<34> sl<54> vdd vss wl<34> / cell_PIM
XI24547 bl<62> cbl<31> in1<16> in2<16> sl<62> vdd vss wl<16> / cell_PIM
XI24546 bl<62> cbl<31> in1<17> in2<17> sl<62> vdd vss wl<17> / cell_PIM
XI24545 bl<62> cbl<31> in1<15> in2<15> sl<62> vdd vss wl<15> / cell_PIM
XI22723 bl<62> cbl<31> in1<73> in2<73> sl<62> vdd vss wl<73> / cell_PIM
XI23273 bl<50> cbl<25> in1<51> in2<51> sl<50> vdd vss wl<51> / cell_PIM
XI23891 bl<52> cbl<26> in1<33> in2<33> sl<52> vdd vss wl<33> / cell_PIM
XI23890 bl<52> cbl<26> in1<32> in2<32> sl<52> vdd vss wl<32> / cell_PIM
XI23889 bl<52> cbl<26> in1<36> in2<36> sl<52> vdd vss wl<36> / cell_PIM
XI24539 bl<60> cbl<30> in1<14> in2<14> sl<60> vdd vss wl<14> / cell_PIM
XI24537 bl<60> cbl<30> in1<17> in2<17> sl<60> vdd vss wl<17> / cell_PIM
XI24536 bl<60> cbl<30> in1<16> in2<16> sl<60> vdd vss wl<16> / cell_PIM
XI24535 bl<60> cbl<30> in1<15> in2<15> sl<60> vdd vss wl<15> / cell_PIM
XI23888 bl<52> cbl<26> in1<35> in2<35> sl<52> vdd vss wl<35> / cell_PIM
XI23887 bl<52> cbl<26> in1<34> in2<34> sl<52> vdd vss wl<34> / cell_PIM
XI23272 bl<50> cbl<25> in1<52> in2<52> sl<50> vdd vss wl<52> / cell_PIM
XI23271 bl<50> cbl<25> in1<54> in2<54> sl<50> vdd vss wl<54> / cell_PIM
XI23270 bl<50> cbl<25> in1<55> in2<55> sl<50> vdd vss wl<55> / cell_PIM
XI23269 bl<50> cbl<25> in1<53> in2<53> sl<50> vdd vss wl<53> / cell_PIM
XI22713 bl<60> cbl<30> in1<74> in2<74> sl<60> vdd vss wl<74> / cell_PIM
XI23881 bl<50> cbl<25> in1<32> in2<32> sl<50> vdd vss wl<32> / cell_PIM
XI23880 bl<50> cbl<25> in1<33> in2<33> sl<50> vdd vss wl<33> / cell_PIM
XI23879 bl<50> cbl<25> in1<35> in2<35> sl<50> vdd vss wl<35> / cell_PIM
XI24529 bl<58> cbl<29> in1<13> in2<13> sl<58> vdd vss wl<13> / cell_PIM
XI23263 bl<48> cbl<24> in1<52> in2<52> sl<48> vdd vss wl<52> / cell_PIM
XI23262 bl<48> cbl<24> in1<51> in2<51> sl<48> vdd vss wl<51> / cell_PIM
XI23261 bl<48> cbl<24> in1<55> in2<55> sl<48> vdd vss wl<55> / cell_PIM
XI23878 bl<50> cbl<25> in1<36> in2<36> sl<50> vdd vss wl<36> / cell_PIM
XI23877 bl<50> cbl<25> in1<34> in2<34> sl<50> vdd vss wl<34> / cell_PIM
XI24527 bl<58> cbl<29> in1<16> in2<16> sl<58> vdd vss wl<16> / cell_PIM
XI24526 bl<58> cbl<29> in1<17> in2<17> sl<58> vdd vss wl<17> / cell_PIM
XI24525 bl<58> cbl<29> in1<15> in2<15> sl<58> vdd vss wl<15> / cell_PIM
XI22703 bl<58> cbl<29> in1<73> in2<73> sl<58> vdd vss wl<73> / cell_PIM
XI23260 bl<48> cbl<24> in1<54> in2<54> sl<48> vdd vss wl<54> / cell_PIM
XI23259 bl<48> cbl<24> in1<53> in2<53> sl<48> vdd vss wl<53> / cell_PIM
XI23871 bl<48> cbl<24> in1<33> in2<33> sl<48> vdd vss wl<33> / cell_PIM
XI23870 bl<48> cbl<24> in1<32> in2<32> sl<48> vdd vss wl<32> / cell_PIM
XI23869 bl<48> cbl<24> in1<36> in2<36> sl<48> vdd vss wl<36> / cell_PIM
XI24519 bl<56> cbl<28> in1<13> in2<13> sl<56> vdd vss wl<13> / cell_PIM
XI24517 bl<56> cbl<28> in1<16> in2<16> sl<56> vdd vss wl<16> / cell_PIM
XI24516 bl<56> cbl<28> in1<17> in2<17> sl<56> vdd vss wl<17> / cell_PIM
XI24515 bl<56> cbl<28> in1<15> in2<15> sl<56> vdd vss wl<15> / cell_PIM
XI23868 bl<48> cbl<24> in1<35> in2<35> sl<48> vdd vss wl<35> / cell_PIM
XI23867 bl<48> cbl<24> in1<34> in2<34> sl<48> vdd vss wl<34> / cell_PIM
XI23253 bl<46> cbl<23> in1<51> in2<51> sl<46> vdd vss wl<51> / cell_PIM
XI22693 bl<56> cbl<28> in1<73> in2<73> sl<56> vdd vss wl<73> / cell_PIM
XI23252 bl<46> cbl<23> in1<52> in2<52> sl<46> vdd vss wl<52> / cell_PIM
XI23251 bl<46> cbl<23> in1<54> in2<54> sl<46> vdd vss wl<54> / cell_PIM
XI23250 bl<46> cbl<23> in1<55> in2<55> sl<46> vdd vss wl<55> / cell_PIM
XI23249 bl<46> cbl<23> in1<53> in2<53> sl<46> vdd vss wl<53> / cell_PIM
XI23861 bl<46> cbl<23> in1<32> in2<32> sl<46> vdd vss wl<32> / cell_PIM
XI23860 bl<46> cbl<23> in1<33> in2<33> sl<46> vdd vss wl<33> / cell_PIM
XI23859 bl<46> cbl<23> in1<35> in2<35> sl<46> vdd vss wl<35> / cell_PIM
XI24509 bl<54> cbl<27> in1<13> in2<13> sl<54> vdd vss wl<13> / cell_PIM
XI23858 bl<46> cbl<23> in1<36> in2<36> sl<46> vdd vss wl<36> / cell_PIM
XI23857 bl<46> cbl<23> in1<34> in2<34> sl<46> vdd vss wl<34> / cell_PIM
XI24507 bl<54> cbl<27> in1<16> in2<16> sl<54> vdd vss wl<16> / cell_PIM
XI24506 bl<54> cbl<27> in1<17> in2<17> sl<54> vdd vss wl<17> / cell_PIM
XI24505 bl<54> cbl<27> in1<15> in2<15> sl<54> vdd vss wl<15> / cell_PIM
XI22683 bl<54> cbl<27> in1<73> in2<73> sl<54> vdd vss wl<73> / cell_PIM
XI23243 bl<44> cbl<22> in1<52> in2<52> sl<44> vdd vss wl<52> / cell_PIM
XI23242 bl<44> cbl<22> in1<51> in2<51> sl<44> vdd vss wl<51> / cell_PIM
XI23241 bl<44> cbl<22> in1<55> in2<55> sl<44> vdd vss wl<55> / cell_PIM
XI23851 bl<44> cbl<22> in1<33> in2<33> sl<44> vdd vss wl<33> / cell_PIM
XI23850 bl<44> cbl<22> in1<32> in2<32> sl<44> vdd vss wl<32> / cell_PIM
XI23849 bl<44> cbl<22> in1<36> in2<36> sl<44> vdd vss wl<36> / cell_PIM
XI24499 bl<52> cbl<26> in1<14> in2<14> sl<52> vdd vss wl<14> / cell_PIM
XI24497 bl<52> cbl<26> in1<17> in2<17> sl<52> vdd vss wl<17> / cell_PIM
XI24496 bl<52> cbl<26> in1<16> in2<16> sl<52> vdd vss wl<16> / cell_PIM
XI24495 bl<52> cbl<26> in1<15> in2<15> sl<52> vdd vss wl<15> / cell_PIM
XI23848 bl<44> cbl<22> in1<35> in2<35> sl<44> vdd vss wl<35> / cell_PIM
XI23847 bl<44> cbl<22> in1<34> in2<34> sl<44> vdd vss wl<34> / cell_PIM
XI23240 bl<44> cbl<22> in1<54> in2<54> sl<44> vdd vss wl<54> / cell_PIM
XI23239 bl<44> cbl<22> in1<53> in2<53> sl<44> vdd vss wl<53> / cell_PIM
XI22673 bl<52> cbl<26> in1<74> in2<74> sl<52> vdd vss wl<74> / cell_PIM
XI23233 bl<42> cbl<21> in1<51> in2<51> sl<42> vdd vss wl<51> / cell_PIM
XI23841 bl<42> cbl<21> in1<32> in2<32> sl<42> vdd vss wl<32> / cell_PIM
XI23840 bl<42> cbl<21> in1<33> in2<33> sl<42> vdd vss wl<33> / cell_PIM
XI23839 bl<42> cbl<21> in1<35> in2<35> sl<42> vdd vss wl<35> / cell_PIM
XI24489 bl<50> cbl<25> in1<13> in2<13> sl<50> vdd vss wl<13> / cell_PIM
XI23232 bl<42> cbl<21> in1<52> in2<52> sl<42> vdd vss wl<52> / cell_PIM
XI23231 bl<42> cbl<21> in1<54> in2<54> sl<42> vdd vss wl<54> / cell_PIM
XI23230 bl<42> cbl<21> in1<55> in2<55> sl<42> vdd vss wl<55> / cell_PIM
XI23229 bl<42> cbl<21> in1<53> in2<53> sl<42> vdd vss wl<53> / cell_PIM
XI23838 bl<42> cbl<21> in1<36> in2<36> sl<42> vdd vss wl<36> / cell_PIM
XI23837 bl<42> cbl<21> in1<34> in2<34> sl<42> vdd vss wl<34> / cell_PIM
XI24487 bl<50> cbl<25> in1<16> in2<16> sl<50> vdd vss wl<16> / cell_PIM
XI24486 bl<50> cbl<25> in1<17> in2<17> sl<50> vdd vss wl<17> / cell_PIM
XI24485 bl<50> cbl<25> in1<15> in2<15> sl<50> vdd vss wl<15> / cell_PIM
XI22663 bl<50> cbl<25> in1<73> in2<73> sl<50> vdd vss wl<73> / cell_PIM
XI23831 bl<40> cbl<20> in1<32> in2<32> sl<40> vdd vss wl<32> / cell_PIM
XI23830 bl<40> cbl<20> in1<33> in2<33> sl<40> vdd vss wl<33> / cell_PIM
XI23829 bl<40> cbl<20> in1<35> in2<35> sl<40> vdd vss wl<35> / cell_PIM
XI24479 bl<48> cbl<24> in1<14> in2<14> sl<48> vdd vss wl<14> / cell_PIM
XI24477 bl<48> cbl<24> in1<17> in2<17> sl<48> vdd vss wl<17> / cell_PIM
XI24476 bl<48> cbl<24> in1<16> in2<16> sl<48> vdd vss wl<16> / cell_PIM
XI24475 bl<48> cbl<24> in1<15> in2<15> sl<48> vdd vss wl<15> / cell_PIM
XI23828 bl<40> cbl<20> in1<36> in2<36> sl<40> vdd vss wl<36> / cell_PIM
XI23827 bl<40> cbl<20> in1<34> in2<34> sl<40> vdd vss wl<34> / cell_PIM
XI23223 bl<40> cbl<20> in1<51> in2<51> sl<40> vdd vss wl<51> / cell_PIM
XI23222 bl<40> cbl<20> in1<52> in2<52> sl<40> vdd vss wl<52> / cell_PIM
XI23221 bl<40> cbl<20> in1<54> in2<54> sl<40> vdd vss wl<54> / cell_PIM
XI22653 bl<48> cbl<24> in1<74> in2<74> sl<48> vdd vss wl<74> / cell_PIM
XI23220 bl<40> cbl<20> in1<55> in2<55> sl<40> vdd vss wl<55> / cell_PIM
XI23219 bl<40> cbl<20> in1<53> in2<53> sl<40> vdd vss wl<53> / cell_PIM
XI23821 bl<38> cbl<19> in1<32> in2<32> sl<38> vdd vss wl<32> / cell_PIM
XI23820 bl<38> cbl<19> in1<33> in2<33> sl<38> vdd vss wl<33> / cell_PIM
XI23819 bl<38> cbl<19> in1<35> in2<35> sl<38> vdd vss wl<35> / cell_PIM
XI24469 bl<46> cbl<23> in1<13> in2<13> sl<46> vdd vss wl<13> / cell_PIM
XI23213 bl<38> cbl<19> in1<51> in2<51> sl<38> vdd vss wl<51> / cell_PIM
XI23818 bl<38> cbl<19> in1<36> in2<36> sl<38> vdd vss wl<36> / cell_PIM
XI23817 bl<38> cbl<19> in1<34> in2<34> sl<38> vdd vss wl<34> / cell_PIM
XI24467 bl<46> cbl<23> in1<16> in2<16> sl<46> vdd vss wl<16> / cell_PIM
XI24466 bl<46> cbl<23> in1<17> in2<17> sl<46> vdd vss wl<17> / cell_PIM
XI24465 bl<46> cbl<23> in1<15> in2<15> sl<46> vdd vss wl<15> / cell_PIM
XI22643 bl<46> cbl<23> in1<73> in2<73> sl<46> vdd vss wl<73> / cell_PIM
XI23212 bl<38> cbl<19> in1<52> in2<52> sl<38> vdd vss wl<52> / cell_PIM
XI23211 bl<38> cbl<19> in1<54> in2<54> sl<38> vdd vss wl<54> / cell_PIM
XI23210 bl<38> cbl<19> in1<55> in2<55> sl<38> vdd vss wl<55> / cell_PIM
XI23209 bl<38> cbl<19> in1<53> in2<53> sl<38> vdd vss wl<53> / cell_PIM
XI23811 bl<36> cbl<18> in1<33> in2<33> sl<36> vdd vss wl<33> / cell_PIM
XI23810 bl<36> cbl<18> in1<32> in2<32> sl<36> vdd vss wl<32> / cell_PIM
XI23809 bl<36> cbl<18> in1<36> in2<36> sl<36> vdd vss wl<36> / cell_PIM
XI24459 bl<44> cbl<22> in1<14> in2<14> sl<44> vdd vss wl<14> / cell_PIM
XI24457 bl<44> cbl<22> in1<17> in2<17> sl<44> vdd vss wl<17> / cell_PIM
XI24456 bl<44> cbl<22> in1<16> in2<16> sl<44> vdd vss wl<16> / cell_PIM
XI24455 bl<44> cbl<22> in1<15> in2<15> sl<44> vdd vss wl<15> / cell_PIM
XI23808 bl<36> cbl<18> in1<35> in2<35> sl<36> vdd vss wl<35> / cell_PIM
XI23807 bl<36> cbl<18> in1<34> in2<34> sl<36> vdd vss wl<34> / cell_PIM
XI22633 bl<44> cbl<22> in1<74> in2<74> sl<44> vdd vss wl<74> / cell_PIM
XI23203 bl<36> cbl<18> in1<52> in2<52> sl<36> vdd vss wl<52> / cell_PIM
XI23202 bl<36> cbl<18> in1<51> in2<51> sl<36> vdd vss wl<51> / cell_PIM
XI23201 bl<36> cbl<18> in1<55> in2<55> sl<36> vdd vss wl<55> / cell_PIM
XI23801 bl<34> cbl<17> in1<32> in2<32> sl<34> vdd vss wl<32> / cell_PIM
XI23800 bl<34> cbl<17> in1<33> in2<33> sl<34> vdd vss wl<33> / cell_PIM
XI23799 bl<34> cbl<17> in1<35> in2<35> sl<34> vdd vss wl<35> / cell_PIM
XI24449 bl<42> cbl<21> in1<13> in2<13> sl<42> vdd vss wl<13> / cell_PIM
XI23200 bl<36> cbl<18> in1<54> in2<54> sl<36> vdd vss wl<54> / cell_PIM
XI23199 bl<36> cbl<18> in1<53> in2<53> sl<36> vdd vss wl<53> / cell_PIM
XI23798 bl<34> cbl<17> in1<36> in2<36> sl<34> vdd vss wl<36> / cell_PIM
XI23797 bl<34> cbl<17> in1<34> in2<34> sl<34> vdd vss wl<34> / cell_PIM
XI24447 bl<42> cbl<21> in1<16> in2<16> sl<42> vdd vss wl<16> / cell_PIM
XI24446 bl<42> cbl<21> in1<17> in2<17> sl<42> vdd vss wl<17> / cell_PIM
XI24445 bl<42> cbl<21> in1<15> in2<15> sl<42> vdd vss wl<15> / cell_PIM
XI22623 bl<42> cbl<21> in1<73> in2<73> sl<42> vdd vss wl<73> / cell_PIM
XI23193 bl<34> cbl<17> in1<51> in2<51> sl<34> vdd vss wl<51> / cell_PIM
XI23791 bl<32> cbl<16> in1<33> in2<33> sl<32> vdd vss wl<33> / cell_PIM
XI23790 bl<32> cbl<16> in1<32> in2<32> sl<32> vdd vss wl<32> / cell_PIM
XI23789 bl<32> cbl<16> in1<36> in2<36> sl<32> vdd vss wl<36> / cell_PIM
XI24439 bl<40> cbl<20> in1<13> in2<13> sl<40> vdd vss wl<13> / cell_PIM
XI24437 bl<40> cbl<20> in1<16> in2<16> sl<40> vdd vss wl<16> / cell_PIM
XI24436 bl<40> cbl<20> in1<17> in2<17> sl<40> vdd vss wl<17> / cell_PIM
XI24435 bl<40> cbl<20> in1<15> in2<15> sl<40> vdd vss wl<15> / cell_PIM
XI23788 bl<32> cbl<16> in1<35> in2<35> sl<32> vdd vss wl<35> / cell_PIM
XI23787 bl<32> cbl<16> in1<34> in2<34> sl<32> vdd vss wl<34> / cell_PIM
XI23192 bl<34> cbl<17> in1<52> in2<52> sl<34> vdd vss wl<52> / cell_PIM
XI23191 bl<34> cbl<17> in1<54> in2<54> sl<34> vdd vss wl<54> / cell_PIM
XI23190 bl<34> cbl<17> in1<55> in2<55> sl<34> vdd vss wl<55> / cell_PIM
XI23189 bl<34> cbl<17> in1<53> in2<53> sl<34> vdd vss wl<53> / cell_PIM
XI22613 bl<40> cbl<20> in1<73> in2<73> sl<40> vdd vss wl<73> / cell_PIM
XI23782 bl<62> cbl<31> in1<37> in2<37> sl<62> vdd vss wl<37> / cell_PIM
XI23781 bl<62> cbl<31> in1<38> in2<38> sl<62> vdd vss wl<38> / cell_PIM
XI23780 bl<62> cbl<31> in1<40> in2<40> sl<62> vdd vss wl<40> / cell_PIM
XI23779 bl<62> cbl<31> in1<39> in2<39> sl<62> vdd vss wl<39> / cell_PIM
XI24429 bl<38> cbl<19> in1<13> in2<13> sl<38> vdd vss wl<13> / cell_PIM
XI23183 bl<32> cbl<16> in1<52> in2<52> sl<32> vdd vss wl<52> / cell_PIM
XI23182 bl<32> cbl<16> in1<51> in2<51> sl<32> vdd vss wl<51> / cell_PIM
XI23181 bl<32> cbl<16> in1<55> in2<55> sl<32> vdd vss wl<55> / cell_PIM
XI23774 bl<60> cbl<30> in1<38> in2<38> sl<60> vdd vss wl<38> / cell_PIM
XI24427 bl<38> cbl<19> in1<16> in2<16> sl<38> vdd vss wl<16> / cell_PIM
XI24426 bl<38> cbl<19> in1<17> in2<17> sl<38> vdd vss wl<17> / cell_PIM
XI24425 bl<38> cbl<19> in1<15> in2<15> sl<38> vdd vss wl<15> / cell_PIM
XI22603 bl<38> cbl<19> in1<73> in2<73> sl<38> vdd vss wl<73> / cell_PIM
XI23180 bl<32> cbl<16> in1<54> in2<54> sl<32> vdd vss wl<54> / cell_PIM
XI23179 bl<32> cbl<16> in1<53> in2<53> sl<32> vdd vss wl<53> / cell_PIM
XI23773 bl<60> cbl<30> in1<37> in2<37> sl<60> vdd vss wl<37> / cell_PIM
XI23772 bl<60> cbl<30> in1<40> in2<40> sl<60> vdd vss wl<40> / cell_PIM
XI23771 bl<60> cbl<30> in1<39> in2<39> sl<60> vdd vss wl<39> / cell_PIM
XI24419 bl<36> cbl<18> in1<14> in2<14> sl<36> vdd vss wl<14> / cell_PIM
XI24417 bl<36> cbl<18> in1<17> in2<17> sl<36> vdd vss wl<17> / cell_PIM
XI24416 bl<36> cbl<18> in1<16> in2<16> sl<36> vdd vss wl<16> / cell_PIM
XI24415 bl<36> cbl<18> in1<15> in2<15> sl<36> vdd vss wl<15> / cell_PIM
XI23766 bl<58> cbl<29> in1<37> in2<37> sl<58> vdd vss wl<37> / cell_PIM
XI23765 bl<58> cbl<29> in1<38> in2<38> sl<58> vdd vss wl<38> / cell_PIM
XI23764 bl<58> cbl<29> in1<40> in2<40> sl<58> vdd vss wl<40> / cell_PIM
XI23173 bl<62> cbl<31> in1<56> in2<56> sl<62> vdd vss wl<56> / cell_PIM
XI22593 bl<36> cbl<18> in1<74> in2<74> sl<36> vdd vss wl<74> / cell_PIM
XI23172 bl<62> cbl<31> in1<57> in2<57> sl<62> vdd vss wl<57> / cell_PIM
XI23171 bl<62> cbl<31> in1<59> in2<59> sl<62> vdd vss wl<59> / cell_PIM
XI23170 bl<62> cbl<31> in1<60> in2<60> sl<62> vdd vss wl<60> / cell_PIM
XI23169 bl<62> cbl<31> in1<58> in2<58> sl<62> vdd vss wl<58> / cell_PIM
XI23763 bl<58> cbl<29> in1<39> in2<39> sl<58> vdd vss wl<39> / cell_PIM
XI24409 bl<34> cbl<17> in1<13> in2<13> sl<34> vdd vss wl<13> / cell_PIM
XI23758 bl<56> cbl<28> in1<37> in2<37> sl<56> vdd vss wl<37> / cell_PIM
XI23757 bl<56> cbl<28> in1<38> in2<38> sl<56> vdd vss wl<38> / cell_PIM
XI23756 bl<56> cbl<28> in1<40> in2<40> sl<56> vdd vss wl<40> / cell_PIM
XI23755 bl<56> cbl<28> in1<39> in2<39> sl<56> vdd vss wl<39> / cell_PIM
XI24407 bl<34> cbl<17> in1<16> in2<16> sl<34> vdd vss wl<16> / cell_PIM
XI24406 bl<34> cbl<17> in1<17> in2<17> sl<34> vdd vss wl<17> / cell_PIM
XI24405 bl<34> cbl<17> in1<15> in2<15> sl<34> vdd vss wl<15> / cell_PIM
XI22583 bl<34> cbl<17> in1<73> in2<73> sl<34> vdd vss wl<73> / cell_PIM
XI23163 bl<60> cbl<30> in1<57> in2<57> sl<60> vdd vss wl<57> / cell_PIM
XI23162 bl<60> cbl<30> in1<56> in2<56> sl<60> vdd vss wl<56> / cell_PIM
XI23161 bl<60> cbl<30> in1<60> in2<60> sl<60> vdd vss wl<60> / cell_PIM
XI23750 bl<54> cbl<27> in1<37> in2<37> sl<54> vdd vss wl<37> / cell_PIM
XI23749 bl<54> cbl<27> in1<38> in2<38> sl<54> vdd vss wl<38> / cell_PIM
XI24399 bl<32> cbl<16> in1<14> in2<14> sl<32> vdd vss wl<14> / cell_PIM
XI24397 bl<32> cbl<16> in1<17> in2<17> sl<32> vdd vss wl<17> / cell_PIM
XI24396 bl<32> cbl<16> in1<16> in2<16> sl<32> vdd vss wl<16> / cell_PIM
XI24395 bl<32> cbl<16> in1<15> in2<15> sl<32> vdd vss wl<15> / cell_PIM
XI23748 bl<54> cbl<27> in1<40> in2<40> sl<54> vdd vss wl<40> / cell_PIM
XI23747 bl<54> cbl<27> in1<39> in2<39> sl<54> vdd vss wl<39> / cell_PIM
XI23160 bl<60> cbl<30> in1<59> in2<59> sl<60> vdd vss wl<59> / cell_PIM
XI23159 bl<60> cbl<30> in1<58> in2<58> sl<60> vdd vss wl<58> / cell_PIM
XI22573 bl<32> cbl<16> in1<74> in2<74> sl<32> vdd vss wl<74> / cell_PIM
XI23153 bl<58> cbl<29> in1<56> in2<56> sl<58> vdd vss wl<56> / cell_PIM
XI23742 bl<52> cbl<26> in1<38> in2<38> sl<52> vdd vss wl<38> / cell_PIM
XI23741 bl<52> cbl<26> in1<37> in2<37> sl<52> vdd vss wl<37> / cell_PIM
XI23740 bl<52> cbl<26> in1<40> in2<40> sl<52> vdd vss wl<40> / cell_PIM
XI23739 bl<52> cbl<26> in1<39> in2<39> sl<52> vdd vss wl<39> / cell_PIM
XI24390 bl<62> cbl<31> in1<18> in2<18> sl<62> vdd vss wl<18> / cell_PIM
XI24389 bl<62> cbl<31> in1<19> in2<19> sl<62> vdd vss wl<19> / cell_PIM
XI23152 bl<58> cbl<29> in1<57> in2<57> sl<58> vdd vss wl<57> / cell_PIM
XI23151 bl<58> cbl<29> in1<59> in2<59> sl<58> vdd vss wl<59> / cell_PIM
XI23150 bl<58> cbl<29> in1<60> in2<60> sl<58> vdd vss wl<60> / cell_PIM
XI23149 bl<58> cbl<29> in1<58> in2<58> sl<58> vdd vss wl<58> / cell_PIM
XI23734 bl<50> cbl<25> in1<37> in2<37> sl<50> vdd vss wl<37> / cell_PIM
XI24387 bl<62> cbl<31> in1<20> in2<20> sl<62> vdd vss wl<20> / cell_PIM
XI21582 bl<48> cbl<24> in1<105> in2<105> sl<48> vdd vss wl<105> / cell_PIM
XI21581 bl<48> cbl<24> in1<104> in2<104> sl<48> vdd vss wl<104> / cell_PIM
XI21580 bl<48> cbl<24> in1<107> in2<107> sl<48> vdd vss wl<107> / cell_PIM
XI21579 bl<48> cbl<24> in1<106> in2<106> sl<48> vdd vss wl<106> / cell_PIM
XI22233 bl<54> cbl<27> in1<87> in2<87> sl<54> vdd vss wl<87> / cell_PIM
XI22882 bl<62> cbl<31> in1<69> in2<69> sl<62> vdd vss wl<69> / cell_PIM
XI22881 bl<62> cbl<31> in1<68> in2<68> sl<62> vdd vss wl<68> / cell_PIM
XI22875 bl<60> cbl<30> in1<67> in2<67> sl<60> vdd vss wl<67> / cell_PIM
XI22227 bl<52> cbl<26> in1<86> in2<86> sl<52> vdd vss wl<86> / cell_PIM
XI22226 bl<52> cbl<26> in1<85> in2<85> sl<52> vdd vss wl<85> / cell_PIM
XI22225 bl<52> cbl<26> in1<84> in2<84> sl<52> vdd vss wl<84> / cell_PIM
XI22224 bl<52> cbl<26> in1<88> in2<88> sl<52> vdd vss wl<88> / cell_PIM
XI21574 bl<46> cbl<23> in1<104> in2<104> sl<46> vdd vss wl<104> / cell_PIM
XI22874 bl<60> cbl<30> in1<66> in2<66> sl<60> vdd vss wl<66> / cell_PIM
XI21573 bl<46> cbl<23> in1<105> in2<105> sl<46> vdd vss wl<105> / cell_PIM
XI21572 bl<46> cbl<23> in1<107> in2<107> sl<46> vdd vss wl<107> / cell_PIM
XI21571 bl<46> cbl<23> in1<106> in2<106> sl<46> vdd vss wl<106> / cell_PIM
XI22223 bl<52> cbl<26> in1<87> in2<87> sl<52> vdd vss wl<87> / cell_PIM
XI22872 bl<60> cbl<30> in1<69> in2<69> sl<60> vdd vss wl<69> / cell_PIM
XI22871 bl<60> cbl<30> in1<68> in2<68> sl<60> vdd vss wl<68> / cell_PIM
XI21566 bl<44> cbl<22> in1<105> in2<105> sl<44> vdd vss wl<105> / cell_PIM
XI21565 bl<44> cbl<22> in1<104> in2<104> sl<44> vdd vss wl<104> / cell_PIM
XI21564 bl<44> cbl<22> in1<107> in2<107> sl<44> vdd vss wl<107> / cell_PIM
XI22217 bl<50> cbl<25> in1<84> in2<84> sl<50> vdd vss wl<84> / cell_PIM
XI22216 bl<50> cbl<25> in1<85> in2<85> sl<50> vdd vss wl<85> / cell_PIM
XI22215 bl<50> cbl<25> in1<86> in2<86> sl<50> vdd vss wl<86> / cell_PIM
XI22214 bl<50> cbl<25> in1<88> in2<88> sl<50> vdd vss wl<88> / cell_PIM
XI22865 bl<58> cbl<29> in1<65> in2<65> sl<58> vdd vss wl<65> / cell_PIM
XI22864 bl<58> cbl<29> in1<66> in2<66> sl<58> vdd vss wl<66> / cell_PIM
XI21563 bl<44> cbl<22> in1<106> in2<106> sl<44> vdd vss wl<106> / cell_PIM
XI22213 bl<50> cbl<25> in1<87> in2<87> sl<50> vdd vss wl<87> / cell_PIM
XI22862 bl<58> cbl<29> in1<69> in2<69> sl<58> vdd vss wl<69> / cell_PIM
XI22861 bl<58> cbl<29> in1<68> in2<68> sl<58> vdd vss wl<68> / cell_PIM
XI22855 bl<56> cbl<28> in1<65> in2<65> sl<56> vdd vss wl<65> / cell_PIM
XI22207 bl<48> cbl<24> in1<86> in2<86> sl<48> vdd vss wl<86> / cell_PIM
XI22206 bl<48> cbl<24> in1<85> in2<85> sl<48> vdd vss wl<85> / cell_PIM
XI22205 bl<48> cbl<24> in1<84> in2<84> sl<48> vdd vss wl<84> / cell_PIM
XI22204 bl<48> cbl<24> in1<88> in2<88> sl<48> vdd vss wl<88> / cell_PIM
XI21558 bl<42> cbl<21> in1<104> in2<104> sl<42> vdd vss wl<104> / cell_PIM
XI21557 bl<42> cbl<21> in1<105> in2<105> sl<42> vdd vss wl<105> / cell_PIM
XI21556 bl<42> cbl<21> in1<107> in2<107> sl<42> vdd vss wl<107> / cell_PIM
XI21555 bl<42> cbl<21> in1<106> in2<106> sl<42> vdd vss wl<106> / cell_PIM
XI22854 bl<56> cbl<28> in1<66> in2<66> sl<56> vdd vss wl<66> / cell_PIM
XI21550 bl<40> cbl<20> in1<104> in2<104> sl<40> vdd vss wl<104> / cell_PIM
XI21549 bl<40> cbl<20> in1<105> in2<105> sl<40> vdd vss wl<105> / cell_PIM
XI22203 bl<48> cbl<24> in1<87> in2<87> sl<48> vdd vss wl<87> / cell_PIM
XI22852 bl<56> cbl<28> in1<69> in2<69> sl<56> vdd vss wl<69> / cell_PIM
XI22851 bl<56> cbl<28> in1<68> in2<68> sl<56> vdd vss wl<68> / cell_PIM
XI21548 bl<40> cbl<20> in1<107> in2<107> sl<40> vdd vss wl<107> / cell_PIM
XI21547 bl<40> cbl<20> in1<106> in2<106> sl<40> vdd vss wl<106> / cell_PIM
XI22197 bl<46> cbl<23> in1<84> in2<84> sl<46> vdd vss wl<84> / cell_PIM
XI22196 bl<46> cbl<23> in1<85> in2<85> sl<46> vdd vss wl<85> / cell_PIM
XI22195 bl<46> cbl<23> in1<86> in2<86> sl<46> vdd vss wl<86> / cell_PIM
XI22194 bl<46> cbl<23> in1<88> in2<88> sl<46> vdd vss wl<88> / cell_PIM
XI22845 bl<54> cbl<27> in1<65> in2<65> sl<54> vdd vss wl<65> / cell_PIM
XI22844 bl<54> cbl<27> in1<66> in2<66> sl<54> vdd vss wl<66> / cell_PIM
XI21542 bl<38> cbl<19> in1<104> in2<104> sl<38> vdd vss wl<104> / cell_PIM
XI21541 bl<38> cbl<19> in1<105> in2<105> sl<38> vdd vss wl<105> / cell_PIM
XI21540 bl<38> cbl<19> in1<107> in2<107> sl<38> vdd vss wl<107> / cell_PIM
XI21539 bl<38> cbl<19> in1<106> in2<106> sl<38> vdd vss wl<106> / cell_PIM
XI22193 bl<46> cbl<23> in1<87> in2<87> sl<46> vdd vss wl<87> / cell_PIM
XI22842 bl<54> cbl<27> in1<69> in2<69> sl<54> vdd vss wl<69> / cell_PIM
XI22841 bl<54> cbl<27> in1<68> in2<68> sl<54> vdd vss wl<68> / cell_PIM
XI22835 bl<52> cbl<26> in1<67> in2<67> sl<52> vdd vss wl<67> / cell_PIM
XI22187 bl<44> cbl<22> in1<86> in2<86> sl<44> vdd vss wl<86> / cell_PIM
XI22186 bl<44> cbl<22> in1<85> in2<85> sl<44> vdd vss wl<85> / cell_PIM
XI22185 bl<44> cbl<22> in1<84> in2<84> sl<44> vdd vss wl<84> / cell_PIM
XI22184 bl<44> cbl<22> in1<88> in2<88> sl<44> vdd vss wl<88> / cell_PIM
XI21534 bl<36> cbl<18> in1<105> in2<105> sl<36> vdd vss wl<105> / cell_PIM
XI22834 bl<52> cbl<26> in1<66> in2<66> sl<52> vdd vss wl<66> / cell_PIM
XI21533 bl<36> cbl<18> in1<104> in2<104> sl<36> vdd vss wl<104> / cell_PIM
XI21532 bl<36> cbl<18> in1<107> in2<107> sl<36> vdd vss wl<107> / cell_PIM
XI21531 bl<36> cbl<18> in1<106> in2<106> sl<36> vdd vss wl<106> / cell_PIM
XI22183 bl<44> cbl<22> in1<87> in2<87> sl<44> vdd vss wl<87> / cell_PIM
XI22832 bl<52> cbl<26> in1<69> in2<69> sl<52> vdd vss wl<69> / cell_PIM
XI22831 bl<52> cbl<26> in1<68> in2<68> sl<52> vdd vss wl<68> / cell_PIM
XI21526 bl<34> cbl<17> in1<104> in2<104> sl<34> vdd vss wl<104> / cell_PIM
XI21525 bl<34> cbl<17> in1<105> in2<105> sl<34> vdd vss wl<105> / cell_PIM
XI21524 bl<34> cbl<17> in1<107> in2<107> sl<34> vdd vss wl<107> / cell_PIM
XI22177 bl<42> cbl<21> in1<84> in2<84> sl<42> vdd vss wl<84> / cell_PIM
XI22176 bl<42> cbl<21> in1<85> in2<85> sl<42> vdd vss wl<85> / cell_PIM
XI22175 bl<42> cbl<21> in1<86> in2<86> sl<42> vdd vss wl<86> / cell_PIM
XI22174 bl<42> cbl<21> in1<88> in2<88> sl<42> vdd vss wl<88> / cell_PIM
XI22825 bl<50> cbl<25> in1<65> in2<65> sl<50> vdd vss wl<65> / cell_PIM
XI22824 bl<50> cbl<25> in1<66> in2<66> sl<50> vdd vss wl<66> / cell_PIM
XI21523 bl<34> cbl<17> in1<106> in2<106> sl<34> vdd vss wl<106> / cell_PIM
XI22173 bl<42> cbl<21> in1<87> in2<87> sl<42> vdd vss wl<87> / cell_PIM
XI22822 bl<50> cbl<25> in1<69> in2<69> sl<50> vdd vss wl<69> / cell_PIM
XI22821 bl<50> cbl<25> in1<68> in2<68> sl<50> vdd vss wl<68> / cell_PIM
XI22815 bl<48> cbl<24> in1<67> in2<67> sl<48> vdd vss wl<67> / cell_PIM
XI22167 bl<40> cbl<20> in1<84> in2<84> sl<40> vdd vss wl<84> / cell_PIM
XI22166 bl<40> cbl<20> in1<85> in2<85> sl<40> vdd vss wl<85> / cell_PIM
XI22165 bl<40> cbl<20> in1<86> in2<86> sl<40> vdd vss wl<86> / cell_PIM
XI22164 bl<40> cbl<20> in1<88> in2<88> sl<40> vdd vss wl<88> / cell_PIM
XI21518 bl<32> cbl<16> in1<105> in2<105> sl<32> vdd vss wl<105> / cell_PIM
XI21517 bl<32> cbl<16> in1<104> in2<104> sl<32> vdd vss wl<104> / cell_PIM
XI21516 bl<32> cbl<16> in1<107> in2<107> sl<32> vdd vss wl<107> / cell_PIM
XI21515 bl<32> cbl<16> in1<106> in2<106> sl<32> vdd vss wl<106> / cell_PIM
XI22814 bl<48> cbl<24> in1<66> in2<66> sl<48> vdd vss wl<66> / cell_PIM
XI21509 bl<62> cbl<31> in1<108> in2<108> sl<62> vdd vss wl<108> / cell_PIM
XI22163 bl<40> cbl<20> in1<87> in2<87> sl<40> vdd vss wl<87> / cell_PIM
XI22812 bl<48> cbl<24> in1<69> in2<69> sl<48> vdd vss wl<69> / cell_PIM
XI22811 bl<48> cbl<24> in1<68> in2<68> sl<48> vdd vss wl<68> / cell_PIM
XI21508 bl<62> cbl<31> in1<109> in2<109> sl<62> vdd vss wl<109> / cell_PIM
XI21507 bl<62> cbl<31> in1<110> in2<110> sl<62> vdd vss wl<110> / cell_PIM
XI21506 bl<62> cbl<31> in1<112> in2<112> sl<62> vdd vss wl<112> / cell_PIM
XI21505 bl<62> cbl<31> in1<111> in2<111> sl<62> vdd vss wl<111> / cell_PIM
XI22157 bl<38> cbl<19> in1<84> in2<84> sl<38> vdd vss wl<84> / cell_PIM
XI22156 bl<38> cbl<19> in1<85> in2<85> sl<38> vdd vss wl<85> / cell_PIM
XI22155 bl<38> cbl<19> in1<86> in2<86> sl<38> vdd vss wl<86> / cell_PIM
XI22154 bl<38> cbl<19> in1<88> in2<88> sl<38> vdd vss wl<88> / cell_PIM
XI22805 bl<46> cbl<23> in1<65> in2<65> sl<46> vdd vss wl<65> / cell_PIM
XI22804 bl<46> cbl<23> in1<66> in2<66> sl<46> vdd vss wl<66> / cell_PIM
XI21499 bl<60> cbl<30> in1<110> in2<110> sl<60> vdd vss wl<110> / cell_PIM
XI22153 bl<38> cbl<19> in1<87> in2<87> sl<38> vdd vss wl<87> / cell_PIM
XI22802 bl<46> cbl<23> in1<69> in2<69> sl<46> vdd vss wl<69> / cell_PIM
XI22801 bl<46> cbl<23> in1<68> in2<68> sl<46> vdd vss wl<68> / cell_PIM
XI22795 bl<44> cbl<22> in1<67> in2<67> sl<44> vdd vss wl<67> / cell_PIM
XI22147 bl<36> cbl<18> in1<86> in2<86> sl<36> vdd vss wl<86> / cell_PIM
XI22146 bl<36> cbl<18> in1<85> in2<85> sl<36> vdd vss wl<85> / cell_PIM
XI22145 bl<36> cbl<18> in1<84> in2<84> sl<36> vdd vss wl<84> / cell_PIM
XI22144 bl<36> cbl<18> in1<88> in2<88> sl<36> vdd vss wl<88> / cell_PIM
XI21498 bl<60> cbl<30> in1<109> in2<109> sl<60> vdd vss wl<109> / cell_PIM
XI21497 bl<60> cbl<30> in1<108> in2<108> sl<60> vdd vss wl<108> / cell_PIM
XI21496 bl<60> cbl<30> in1<112> in2<112> sl<60> vdd vss wl<112> / cell_PIM
XI21495 bl<60> cbl<30> in1<111> in2<111> sl<60> vdd vss wl<111> / cell_PIM
XI22794 bl<44> cbl<22> in1<66> in2<66> sl<44> vdd vss wl<66> / cell_PIM
XI21489 bl<58> cbl<29> in1<108> in2<108> sl<58> vdd vss wl<108> / cell_PIM
XI22143 bl<36> cbl<18> in1<87> in2<87> sl<36> vdd vss wl<87> / cell_PIM
XI22792 bl<44> cbl<22> in1<69> in2<69> sl<44> vdd vss wl<69> / cell_PIM
XI22791 bl<44> cbl<22> in1<68> in2<68> sl<44> vdd vss wl<68> / cell_PIM
XI21488 bl<58> cbl<29> in1<109> in2<109> sl<58> vdd vss wl<109> / cell_PIM
XI21487 bl<58> cbl<29> in1<110> in2<110> sl<58> vdd vss wl<110> / cell_PIM
XI21486 bl<58> cbl<29> in1<112> in2<112> sl<58> vdd vss wl<112> / cell_PIM
XI21485 bl<58> cbl<29> in1<111> in2<111> sl<58> vdd vss wl<111> / cell_PIM
XI22137 bl<34> cbl<17> in1<84> in2<84> sl<34> vdd vss wl<84> / cell_PIM
XI22136 bl<34> cbl<17> in1<85> in2<85> sl<34> vdd vss wl<85> / cell_PIM
XI22135 bl<34> cbl<17> in1<86> in2<86> sl<34> vdd vss wl<86> / cell_PIM
XI22134 bl<34> cbl<17> in1<88> in2<88> sl<34> vdd vss wl<88> / cell_PIM
XI22785 bl<42> cbl<21> in1<65> in2<65> sl<42> vdd vss wl<65> / cell_PIM
XI22784 bl<42> cbl<21> in1<66> in2<66> sl<42> vdd vss wl<66> / cell_PIM
XI21479 bl<56> cbl<28> in1<108> in2<108> sl<56> vdd vss wl<108> / cell_PIM
XI22133 bl<34> cbl<17> in1<87> in2<87> sl<34> vdd vss wl<87> / cell_PIM
XI22782 bl<42> cbl<21> in1<69> in2<69> sl<42> vdd vss wl<69> / cell_PIM
XI22781 bl<42> cbl<21> in1<68> in2<68> sl<42> vdd vss wl<68> / cell_PIM
XI22775 bl<40> cbl<20> in1<65> in2<65> sl<40> vdd vss wl<65> / cell_PIM
XI22127 bl<32> cbl<16> in1<86> in2<86> sl<32> vdd vss wl<86> / cell_PIM
XI22126 bl<32> cbl<16> in1<85> in2<85> sl<32> vdd vss wl<85> / cell_PIM
XI22125 bl<32> cbl<16> in1<84> in2<84> sl<32> vdd vss wl<84> / cell_PIM
XI22124 bl<32> cbl<16> in1<88> in2<88> sl<32> vdd vss wl<88> / cell_PIM
XI21478 bl<56> cbl<28> in1<109> in2<109> sl<56> vdd vss wl<109> / cell_PIM
XI21477 bl<56> cbl<28> in1<110> in2<110> sl<56> vdd vss wl<110> / cell_PIM
XI21476 bl<56> cbl<28> in1<112> in2<112> sl<56> vdd vss wl<112> / cell_PIM
XI21475 bl<56> cbl<28> in1<111> in2<111> sl<56> vdd vss wl<111> / cell_PIM
XI22774 bl<40> cbl<20> in1<66> in2<66> sl<40> vdd vss wl<66> / cell_PIM
XI21469 bl<54> cbl<27> in1<108> in2<108> sl<54> vdd vss wl<108> / cell_PIM
XI22123 bl<32> cbl<16> in1<87> in2<87> sl<32> vdd vss wl<87> / cell_PIM
XI22772 bl<40> cbl<20> in1<69> in2<69> sl<40> vdd vss wl<69> / cell_PIM
XI22771 bl<40> cbl<20> in1<68> in2<68> sl<40> vdd vss wl<68> / cell_PIM
XI21468 bl<54> cbl<27> in1<109> in2<109> sl<54> vdd vss wl<109> / cell_PIM
XI21467 bl<54> cbl<27> in1<110> in2<110> sl<54> vdd vss wl<110> / cell_PIM
XI21466 bl<54> cbl<27> in1<112> in2<112> sl<54> vdd vss wl<112> / cell_PIM
XI21465 bl<54> cbl<27> in1<111> in2<111> sl<54> vdd vss wl<111> / cell_PIM
XI22117 bl<62> cbl<31> in1<89> in2<89> sl<62> vdd vss wl<89> / cell_PIM
XI22116 bl<62> cbl<31> in1<90> in2<90> sl<62> vdd vss wl<90> / cell_PIM
XI22115 bl<62> cbl<31> in1<91> in2<91> sl<62> vdd vss wl<91> / cell_PIM
XI22114 bl<62> cbl<31> in1<93> in2<93> sl<62> vdd vss wl<93> / cell_PIM
XI22765 bl<38> cbl<19> in1<65> in2<65> sl<38> vdd vss wl<65> / cell_PIM
XI22764 bl<38> cbl<19> in1<66> in2<66> sl<38> vdd vss wl<66> / cell_PIM
XI21459 bl<52> cbl<26> in1<110> in2<110> sl<52> vdd vss wl<110> / cell_PIM
XI22113 bl<62> cbl<31> in1<92> in2<92> sl<62> vdd vss wl<92> / cell_PIM
XI22762 bl<38> cbl<19> in1<69> in2<69> sl<38> vdd vss wl<69> / cell_PIM
XI22761 bl<38> cbl<19> in1<68> in2<68> sl<38> vdd vss wl<68> / cell_PIM
XI22755 bl<36> cbl<18> in1<67> in2<67> sl<36> vdd vss wl<67> / cell_PIM
XI22107 bl<60> cbl<30> in1<91> in2<91> sl<60> vdd vss wl<91> / cell_PIM
XI22106 bl<60> cbl<30> in1<90> in2<90> sl<60> vdd vss wl<90> / cell_PIM
XI22105 bl<60> cbl<30> in1<89> in2<89> sl<60> vdd vss wl<89> / cell_PIM
XI22104 bl<60> cbl<30> in1<93> in2<93> sl<60> vdd vss wl<93> / cell_PIM
XI21458 bl<52> cbl<26> in1<109> in2<109> sl<52> vdd vss wl<109> / cell_PIM
XI21457 bl<52> cbl<26> in1<108> in2<108> sl<52> vdd vss wl<108> / cell_PIM
XI21456 bl<52> cbl<26> in1<112> in2<112> sl<52> vdd vss wl<112> / cell_PIM
XI21455 bl<52> cbl<26> in1<111> in2<111> sl<52> vdd vss wl<111> / cell_PIM
XI22754 bl<36> cbl<18> in1<66> in2<66> sl<36> vdd vss wl<66> / cell_PIM
XI21449 bl<50> cbl<25> in1<108> in2<108> sl<50> vdd vss wl<108> / cell_PIM
XI22103 bl<60> cbl<30> in1<92> in2<92> sl<60> vdd vss wl<92> / cell_PIM
XI22752 bl<36> cbl<18> in1<69> in2<69> sl<36> vdd vss wl<69> / cell_PIM
XI22751 bl<36> cbl<18> in1<68> in2<68> sl<36> vdd vss wl<68> / cell_PIM
XI21448 bl<50> cbl<25> in1<109> in2<109> sl<50> vdd vss wl<109> / cell_PIM
XI21447 bl<50> cbl<25> in1<110> in2<110> sl<50> vdd vss wl<110> / cell_PIM
XI21446 bl<50> cbl<25> in1<112> in2<112> sl<50> vdd vss wl<112> / cell_PIM
XI21445 bl<50> cbl<25> in1<111> in2<111> sl<50> vdd vss wl<111> / cell_PIM
XI22097 bl<58> cbl<29> in1<89> in2<89> sl<58> vdd vss wl<89> / cell_PIM
XI22096 bl<58> cbl<29> in1<90> in2<90> sl<58> vdd vss wl<90> / cell_PIM
XI22095 bl<58> cbl<29> in1<91> in2<91> sl<58> vdd vss wl<91> / cell_PIM
XI22094 bl<58> cbl<29> in1<93> in2<93> sl<58> vdd vss wl<93> / cell_PIM
XI22745 bl<34> cbl<17> in1<65> in2<65> sl<34> vdd vss wl<65> / cell_PIM
XI22744 bl<34> cbl<17> in1<66> in2<66> sl<34> vdd vss wl<66> / cell_PIM
XI21439 bl<48> cbl<24> in1<110> in2<110> sl<48> vdd vss wl<110> / cell_PIM
XI22093 bl<58> cbl<29> in1<92> in2<92> sl<58> vdd vss wl<92> / cell_PIM
XI22742 bl<34> cbl<17> in1<69> in2<69> sl<34> vdd vss wl<69> / cell_PIM
XI22741 bl<34> cbl<17> in1<68> in2<68> sl<34> vdd vss wl<68> / cell_PIM
XI22735 bl<32> cbl<16> in1<67> in2<67> sl<32> vdd vss wl<67> / cell_PIM
XI22087 bl<56> cbl<28> in1<89> in2<89> sl<56> vdd vss wl<89> / cell_PIM
XI22086 bl<56> cbl<28> in1<90> in2<90> sl<56> vdd vss wl<90> / cell_PIM
XI22085 bl<56> cbl<28> in1<91> in2<91> sl<56> vdd vss wl<91> / cell_PIM
XI22084 bl<56> cbl<28> in1<93> in2<93> sl<56> vdd vss wl<93> / cell_PIM
XI21438 bl<48> cbl<24> in1<109> in2<109> sl<48> vdd vss wl<109> / cell_PIM
XI21437 bl<48> cbl<24> in1<108> in2<108> sl<48> vdd vss wl<108> / cell_PIM
XI21436 bl<48> cbl<24> in1<112> in2<112> sl<48> vdd vss wl<112> / cell_PIM
XI21435 bl<48> cbl<24> in1<111> in2<111> sl<48> vdd vss wl<111> / cell_PIM
XI22734 bl<32> cbl<16> in1<66> in2<66> sl<32> vdd vss wl<66> / cell_PIM
XI21429 bl<46> cbl<23> in1<108> in2<108> sl<46> vdd vss wl<108> / cell_PIM
XI22083 bl<56> cbl<28> in1<92> in2<92> sl<56> vdd vss wl<92> / cell_PIM
XI22732 bl<32> cbl<16> in1<69> in2<69> sl<32> vdd vss wl<69> / cell_PIM
XI22731 bl<32> cbl<16> in1<68> in2<68> sl<32> vdd vss wl<68> / cell_PIM
XI21428 bl<46> cbl<23> in1<109> in2<109> sl<46> vdd vss wl<109> / cell_PIM
XI21427 bl<46> cbl<23> in1<110> in2<110> sl<46> vdd vss wl<110> / cell_PIM
XI21426 bl<46> cbl<23> in1<112> in2<112> sl<46> vdd vss wl<112> / cell_PIM
XI21425 bl<46> cbl<23> in1<111> in2<111> sl<46> vdd vss wl<111> / cell_PIM
XI22077 bl<54> cbl<27> in1<89> in2<89> sl<54> vdd vss wl<89> / cell_PIM
XI22076 bl<54> cbl<27> in1<90> in2<90> sl<54> vdd vss wl<90> / cell_PIM
XI22075 bl<54> cbl<27> in1<91> in2<91> sl<54> vdd vss wl<91> / cell_PIM
XI22074 bl<54> cbl<27> in1<93> in2<93> sl<54> vdd vss wl<93> / cell_PIM
XI22725 bl<62> cbl<31> in1<70> in2<70> sl<62> vdd vss wl<70> / cell_PIM
XI22724 bl<62> cbl<31> in1<71> in2<71> sl<62> vdd vss wl<71> / cell_PIM
XI21419 bl<44> cbl<22> in1<110> in2<110> sl<44> vdd vss wl<110> / cell_PIM
XI22073 bl<54> cbl<27> in1<92> in2<92> sl<54> vdd vss wl<92> / cell_PIM
XI22722 bl<62> cbl<31> in1<74> in2<74> sl<62> vdd vss wl<74> / cell_PIM
XI22721 bl<62> cbl<31> in1<72> in2<72> sl<62> vdd vss wl<72> / cell_PIM
XI22715 bl<60> cbl<30> in1<71> in2<71> sl<60> vdd vss wl<71> / cell_PIM
XI22067 bl<52> cbl<26> in1<91> in2<91> sl<52> vdd vss wl<91> / cell_PIM
XI22066 bl<52> cbl<26> in1<90> in2<90> sl<52> vdd vss wl<90> / cell_PIM
XI22065 bl<52> cbl<26> in1<89> in2<89> sl<52> vdd vss wl<89> / cell_PIM
XI22064 bl<52> cbl<26> in1<93> in2<93> sl<52> vdd vss wl<93> / cell_PIM
XI21418 bl<44> cbl<22> in1<109> in2<109> sl<44> vdd vss wl<109> / cell_PIM
XI21417 bl<44> cbl<22> in1<108> in2<108> sl<44> vdd vss wl<108> / cell_PIM
XI21416 bl<44> cbl<22> in1<112> in2<112> sl<44> vdd vss wl<112> / cell_PIM
XI21415 bl<44> cbl<22> in1<111> in2<111> sl<44> vdd vss wl<111> / cell_PIM
XI22714 bl<60> cbl<30> in1<70> in2<70> sl<60> vdd vss wl<70> / cell_PIM
XI21409 bl<42> cbl<21> in1<108> in2<108> sl<42> vdd vss wl<108> / cell_PIM
XI22063 bl<52> cbl<26> in1<92> in2<92> sl<52> vdd vss wl<92> / cell_PIM
XI22712 bl<60> cbl<30> in1<73> in2<73> sl<60> vdd vss wl<73> / cell_PIM
XI22711 bl<60> cbl<30> in1<72> in2<72> sl<60> vdd vss wl<72> / cell_PIM
XI21408 bl<42> cbl<21> in1<109> in2<109> sl<42> vdd vss wl<109> / cell_PIM
XI21407 bl<42> cbl<21> in1<110> in2<110> sl<42> vdd vss wl<110> / cell_PIM
XI21406 bl<42> cbl<21> in1<112> in2<112> sl<42> vdd vss wl<112> / cell_PIM
XI21405 bl<42> cbl<21> in1<111> in2<111> sl<42> vdd vss wl<111> / cell_PIM
XI22057 bl<50> cbl<25> in1<89> in2<89> sl<50> vdd vss wl<89> / cell_PIM
XI22056 bl<50> cbl<25> in1<90> in2<90> sl<50> vdd vss wl<90> / cell_PIM
XI22055 bl<50> cbl<25> in1<91> in2<91> sl<50> vdd vss wl<91> / cell_PIM
XI22054 bl<50> cbl<25> in1<93> in2<93> sl<50> vdd vss wl<93> / cell_PIM
XI22705 bl<58> cbl<29> in1<70> in2<70> sl<58> vdd vss wl<70> / cell_PIM
XI22704 bl<58> cbl<29> in1<71> in2<71> sl<58> vdd vss wl<71> / cell_PIM
XI21399 bl<40> cbl<20> in1<108> in2<108> sl<40> vdd vss wl<108> / cell_PIM
XI22053 bl<50> cbl<25> in1<92> in2<92> sl<50> vdd vss wl<92> / cell_PIM
XI22702 bl<58> cbl<29> in1<74> in2<74> sl<58> vdd vss wl<74> / cell_PIM
XI22701 bl<58> cbl<29> in1<72> in2<72> sl<58> vdd vss wl<72> / cell_PIM
XI22695 bl<56> cbl<28> in1<70> in2<70> sl<56> vdd vss wl<70> / cell_PIM
XI22047 bl<48> cbl<24> in1<91> in2<91> sl<48> vdd vss wl<91> / cell_PIM
XI22046 bl<48> cbl<24> in1<90> in2<90> sl<48> vdd vss wl<90> / cell_PIM
XI22045 bl<48> cbl<24> in1<89> in2<89> sl<48> vdd vss wl<89> / cell_PIM
XI22044 bl<48> cbl<24> in1<93> in2<93> sl<48> vdd vss wl<93> / cell_PIM
XI21398 bl<40> cbl<20> in1<109> in2<109> sl<40> vdd vss wl<109> / cell_PIM
XI21397 bl<40> cbl<20> in1<110> in2<110> sl<40> vdd vss wl<110> / cell_PIM
XI21396 bl<40> cbl<20> in1<112> in2<112> sl<40> vdd vss wl<112> / cell_PIM
XI21395 bl<40> cbl<20> in1<111> in2<111> sl<40> vdd vss wl<111> / cell_PIM
XI22694 bl<56> cbl<28> in1<71> in2<71> sl<56> vdd vss wl<71> / cell_PIM
XI21389 bl<38> cbl<19> in1<108> in2<108> sl<38> vdd vss wl<108> / cell_PIM
XI22043 bl<48> cbl<24> in1<92> in2<92> sl<48> vdd vss wl<92> / cell_PIM
XI22692 bl<56> cbl<28> in1<74> in2<74> sl<56> vdd vss wl<74> / cell_PIM
XI22691 bl<56> cbl<28> in1<72> in2<72> sl<56> vdd vss wl<72> / cell_PIM
XI21388 bl<38> cbl<19> in1<109> in2<109> sl<38> vdd vss wl<109> / cell_PIM
XI21387 bl<38> cbl<19> in1<110> in2<110> sl<38> vdd vss wl<110> / cell_PIM
XI21386 bl<38> cbl<19> in1<112> in2<112> sl<38> vdd vss wl<112> / cell_PIM
XI21385 bl<38> cbl<19> in1<111> in2<111> sl<38> vdd vss wl<111> / cell_PIM
XI22037 bl<46> cbl<23> in1<89> in2<89> sl<46> vdd vss wl<89> / cell_PIM
XI22036 bl<46> cbl<23> in1<90> in2<90> sl<46> vdd vss wl<90> / cell_PIM
XI22035 bl<46> cbl<23> in1<91> in2<91> sl<46> vdd vss wl<91> / cell_PIM
XI22034 bl<46> cbl<23> in1<93> in2<93> sl<46> vdd vss wl<93> / cell_PIM
XI22685 bl<54> cbl<27> in1<70> in2<70> sl<54> vdd vss wl<70> / cell_PIM
XI22684 bl<54> cbl<27> in1<71> in2<71> sl<54> vdd vss wl<71> / cell_PIM
XI21379 bl<36> cbl<18> in1<110> in2<110> sl<36> vdd vss wl<110> / cell_PIM
XI22033 bl<46> cbl<23> in1<92> in2<92> sl<46> vdd vss wl<92> / cell_PIM
XI22682 bl<54> cbl<27> in1<74> in2<74> sl<54> vdd vss wl<74> / cell_PIM
XI22681 bl<54> cbl<27> in1<72> in2<72> sl<54> vdd vss wl<72> / cell_PIM
XI22675 bl<52> cbl<26> in1<71> in2<71> sl<52> vdd vss wl<71> / cell_PIM
XI22027 bl<44> cbl<22> in1<91> in2<91> sl<44> vdd vss wl<91> / cell_PIM
XI22026 bl<44> cbl<22> in1<90> in2<90> sl<44> vdd vss wl<90> / cell_PIM
XI22025 bl<44> cbl<22> in1<89> in2<89> sl<44> vdd vss wl<89> / cell_PIM
XI22024 bl<44> cbl<22> in1<93> in2<93> sl<44> vdd vss wl<93> / cell_PIM
XI21378 bl<36> cbl<18> in1<109> in2<109> sl<36> vdd vss wl<109> / cell_PIM
XI21377 bl<36> cbl<18> in1<108> in2<108> sl<36> vdd vss wl<108> / cell_PIM
XI21376 bl<36> cbl<18> in1<112> in2<112> sl<36> vdd vss wl<112> / cell_PIM
XI21375 bl<36> cbl<18> in1<111> in2<111> sl<36> vdd vss wl<111> / cell_PIM
XI22674 bl<52> cbl<26> in1<70> in2<70> sl<52> vdd vss wl<70> / cell_PIM
XI21369 bl<34> cbl<17> in1<108> in2<108> sl<34> vdd vss wl<108> / cell_PIM
XI22023 bl<44> cbl<22> in1<92> in2<92> sl<44> vdd vss wl<92> / cell_PIM
XI22672 bl<52> cbl<26> in1<73> in2<73> sl<52> vdd vss wl<73> / cell_PIM
XI22671 bl<52> cbl<26> in1<72> in2<72> sl<52> vdd vss wl<72> / cell_PIM
XI21368 bl<34> cbl<17> in1<109> in2<109> sl<34> vdd vss wl<109> / cell_PIM
XI21367 bl<34> cbl<17> in1<110> in2<110> sl<34> vdd vss wl<110> / cell_PIM
XI21366 bl<34> cbl<17> in1<112> in2<112> sl<34> vdd vss wl<112> / cell_PIM
XI21365 bl<34> cbl<17> in1<111> in2<111> sl<34> vdd vss wl<111> / cell_PIM
XI22017 bl<42> cbl<21> in1<89> in2<89> sl<42> vdd vss wl<89> / cell_PIM
XI22016 bl<42> cbl<21> in1<90> in2<90> sl<42> vdd vss wl<90> / cell_PIM
XI22015 bl<42> cbl<21> in1<91> in2<91> sl<42> vdd vss wl<91> / cell_PIM
XI22014 bl<42> cbl<21> in1<93> in2<93> sl<42> vdd vss wl<93> / cell_PIM
XI22665 bl<50> cbl<25> in1<70> in2<70> sl<50> vdd vss wl<70> / cell_PIM
XI22664 bl<50> cbl<25> in1<71> in2<71> sl<50> vdd vss wl<71> / cell_PIM
XI21359 bl<32> cbl<16> in1<110> in2<110> sl<32> vdd vss wl<110> / cell_PIM
XI22013 bl<42> cbl<21> in1<92> in2<92> sl<42> vdd vss wl<92> / cell_PIM
XI22662 bl<50> cbl<25> in1<74> in2<74> sl<50> vdd vss wl<74> / cell_PIM
XI22661 bl<50> cbl<25> in1<72> in2<72> sl<50> vdd vss wl<72> / cell_PIM
XI22655 bl<48> cbl<24> in1<71> in2<71> sl<48> vdd vss wl<71> / cell_PIM
XI22007 bl<40> cbl<20> in1<89> in2<89> sl<40> vdd vss wl<89> / cell_PIM
XI22006 bl<40> cbl<20> in1<90> in2<90> sl<40> vdd vss wl<90> / cell_PIM
XI22005 bl<40> cbl<20> in1<91> in2<91> sl<40> vdd vss wl<91> / cell_PIM
XI22004 bl<40> cbl<20> in1<93> in2<93> sl<40> vdd vss wl<93> / cell_PIM
XI21358 bl<32> cbl<16> in1<109> in2<109> sl<32> vdd vss wl<109> / cell_PIM
XI21357 bl<32> cbl<16> in1<108> in2<108> sl<32> vdd vss wl<108> / cell_PIM
XI21356 bl<32> cbl<16> in1<112> in2<112> sl<32> vdd vss wl<112> / cell_PIM
XI21355 bl<32> cbl<16> in1<111> in2<111> sl<32> vdd vss wl<111> / cell_PIM
XI22654 bl<48> cbl<24> in1<70> in2<70> sl<48> vdd vss wl<70> / cell_PIM
XI21349 bl<62> cbl<31> in1<113> in2<113> sl<62> vdd vss wl<113> / cell_PIM
XI22003 bl<40> cbl<20> in1<92> in2<92> sl<40> vdd vss wl<92> / cell_PIM
XI22652 bl<48> cbl<24> in1<73> in2<73> sl<48> vdd vss wl<73> / cell_PIM
XI22651 bl<48> cbl<24> in1<72> in2<72> sl<48> vdd vss wl<72> / cell_PIM
XI21348 bl<62> cbl<31> in1<114> in2<114> sl<62> vdd vss wl<114> / cell_PIM
XI21347 bl<62> cbl<31> in1<115> in2<115> sl<62> vdd vss wl<115> / cell_PIM
XI21346 bl<62> cbl<31> in1<117> in2<117> sl<62> vdd vss wl<117> / cell_PIM
XI21345 bl<62> cbl<31> in1<116> in2<116> sl<62> vdd vss wl<116> / cell_PIM
XI21997 bl<38> cbl<19> in1<89> in2<89> sl<38> vdd vss wl<89> / cell_PIM
XI21996 bl<38> cbl<19> in1<90> in2<90> sl<38> vdd vss wl<90> / cell_PIM
XI21995 bl<38> cbl<19> in1<91> in2<91> sl<38> vdd vss wl<91> / cell_PIM
XI21994 bl<38> cbl<19> in1<93> in2<93> sl<38> vdd vss wl<93> / cell_PIM
XI22645 bl<46> cbl<23> in1<70> in2<70> sl<46> vdd vss wl<70> / cell_PIM
XI22644 bl<46> cbl<23> in1<71> in2<71> sl<46> vdd vss wl<71> / cell_PIM
XI21339 bl<60> cbl<30> in1<115> in2<115> sl<60> vdd vss wl<115> / cell_PIM
XI21993 bl<38> cbl<19> in1<92> in2<92> sl<38> vdd vss wl<92> / cell_PIM
XI22642 bl<46> cbl<23> in1<74> in2<74> sl<46> vdd vss wl<74> / cell_PIM
XI22641 bl<46> cbl<23> in1<72> in2<72> sl<46> vdd vss wl<72> / cell_PIM
XI22635 bl<44> cbl<22> in1<71> in2<71> sl<44> vdd vss wl<71> / cell_PIM
XI21987 bl<36> cbl<18> in1<91> in2<91> sl<36> vdd vss wl<91> / cell_PIM
XI21986 bl<36> cbl<18> in1<90> in2<90> sl<36> vdd vss wl<90> / cell_PIM
XI21985 bl<36> cbl<18> in1<89> in2<89> sl<36> vdd vss wl<89> / cell_PIM
XI21984 bl<36> cbl<18> in1<93> in2<93> sl<36> vdd vss wl<93> / cell_PIM
XI21338 bl<60> cbl<30> in1<114> in2<114> sl<60> vdd vss wl<114> / cell_PIM
XI21337 bl<60> cbl<30> in1<113> in2<113> sl<60> vdd vss wl<113> / cell_PIM
XI21336 bl<60> cbl<30> in1<117> in2<117> sl<60> vdd vss wl<117> / cell_PIM
XI21335 bl<60> cbl<30> in1<116> in2<116> sl<60> vdd vss wl<116> / cell_PIM
XI22634 bl<44> cbl<22> in1<70> in2<70> sl<44> vdd vss wl<70> / cell_PIM
XI21329 bl<58> cbl<29> in1<113> in2<113> sl<58> vdd vss wl<113> / cell_PIM
XI21983 bl<36> cbl<18> in1<92> in2<92> sl<36> vdd vss wl<92> / cell_PIM
XI22632 bl<44> cbl<22> in1<73> in2<73> sl<44> vdd vss wl<73> / cell_PIM
XI22631 bl<44> cbl<22> in1<72> in2<72> sl<44> vdd vss wl<72> / cell_PIM
XI21328 bl<58> cbl<29> in1<114> in2<114> sl<58> vdd vss wl<114> / cell_PIM
XI21327 bl<58> cbl<29> in1<115> in2<115> sl<58> vdd vss wl<115> / cell_PIM
XI21326 bl<58> cbl<29> in1<117> in2<117> sl<58> vdd vss wl<117> / cell_PIM
XI21325 bl<58> cbl<29> in1<116> in2<116> sl<58> vdd vss wl<116> / cell_PIM
XI21977 bl<34> cbl<17> in1<89> in2<89> sl<34> vdd vss wl<89> / cell_PIM
XI21976 bl<34> cbl<17> in1<90> in2<90> sl<34> vdd vss wl<90> / cell_PIM
XI21975 bl<34> cbl<17> in1<91> in2<91> sl<34> vdd vss wl<91> / cell_PIM
XI21974 bl<34> cbl<17> in1<93> in2<93> sl<34> vdd vss wl<93> / cell_PIM
XI22625 bl<42> cbl<21> in1<70> in2<70> sl<42> vdd vss wl<70> / cell_PIM
XI22624 bl<42> cbl<21> in1<71> in2<71> sl<42> vdd vss wl<71> / cell_PIM
XI21319 bl<56> cbl<28> in1<113> in2<113> sl<56> vdd vss wl<113> / cell_PIM
XI21973 bl<34> cbl<17> in1<92> in2<92> sl<34> vdd vss wl<92> / cell_PIM
XI22622 bl<42> cbl<21> in1<74> in2<74> sl<42> vdd vss wl<74> / cell_PIM
XI22621 bl<42> cbl<21> in1<72> in2<72> sl<42> vdd vss wl<72> / cell_PIM
XI22615 bl<40> cbl<20> in1<70> in2<70> sl<40> vdd vss wl<70> / cell_PIM
XI21967 bl<32> cbl<16> in1<91> in2<91> sl<32> vdd vss wl<91> / cell_PIM
XI21966 bl<32> cbl<16> in1<90> in2<90> sl<32> vdd vss wl<90> / cell_PIM
XI21965 bl<32> cbl<16> in1<89> in2<89> sl<32> vdd vss wl<89> / cell_PIM
XI21964 bl<32> cbl<16> in1<93> in2<93> sl<32> vdd vss wl<93> / cell_PIM
XI21318 bl<56> cbl<28> in1<114> in2<114> sl<56> vdd vss wl<114> / cell_PIM
XI21317 bl<56> cbl<28> in1<115> in2<115> sl<56> vdd vss wl<115> / cell_PIM
XI21316 bl<56> cbl<28> in1<117> in2<117> sl<56> vdd vss wl<117> / cell_PIM
XI21315 bl<56> cbl<28> in1<116> in2<116> sl<56> vdd vss wl<116> / cell_PIM
XI22614 bl<40> cbl<20> in1<71> in2<71> sl<40> vdd vss wl<71> / cell_PIM
XI21309 bl<54> cbl<27> in1<113> in2<113> sl<54> vdd vss wl<113> / cell_PIM
XI21963 bl<32> cbl<16> in1<92> in2<92> sl<32> vdd vss wl<92> / cell_PIM
XI22612 bl<40> cbl<20> in1<74> in2<74> sl<40> vdd vss wl<74> / cell_PIM
XI22611 bl<40> cbl<20> in1<72> in2<72> sl<40> vdd vss wl<72> / cell_PIM
XI21308 bl<54> cbl<27> in1<114> in2<114> sl<54> vdd vss wl<114> / cell_PIM
XI21307 bl<54> cbl<27> in1<115> in2<115> sl<54> vdd vss wl<115> / cell_PIM
XI21306 bl<54> cbl<27> in1<117> in2<117> sl<54> vdd vss wl<117> / cell_PIM
XI21305 bl<54> cbl<27> in1<116> in2<116> sl<54> vdd vss wl<116> / cell_PIM
XI21957 bl<62> cbl<31> in1<94> in2<94> sl<62> vdd vss wl<94> / cell_PIM
XI21956 bl<62> cbl<31> in1<95> in2<95> sl<62> vdd vss wl<95> / cell_PIM
XI21955 bl<62> cbl<31> in1<97> in2<97> sl<62> vdd vss wl<97> / cell_PIM
XI21954 bl<62> cbl<31> in1<98> in2<98> sl<62> vdd vss wl<98> / cell_PIM
XI22605 bl<38> cbl<19> in1<70> in2<70> sl<38> vdd vss wl<70> / cell_PIM
XI22604 bl<38> cbl<19> in1<71> in2<71> sl<38> vdd vss wl<71> / cell_PIM
XI21299 bl<52> cbl<26> in1<115> in2<115> sl<52> vdd vss wl<115> / cell_PIM
XI21953 bl<62> cbl<31> in1<96> in2<96> sl<62> vdd vss wl<96> / cell_PIM
XI22602 bl<38> cbl<19> in1<74> in2<74> sl<38> vdd vss wl<74> / cell_PIM
XI22601 bl<38> cbl<19> in1<72> in2<72> sl<38> vdd vss wl<72> / cell_PIM
XI22595 bl<36> cbl<18> in1<71> in2<71> sl<36> vdd vss wl<71> / cell_PIM
XI21947 bl<60> cbl<30> in1<95> in2<95> sl<60> vdd vss wl<95> / cell_PIM
XI21946 bl<60> cbl<30> in1<94> in2<94> sl<60> vdd vss wl<94> / cell_PIM
XI21945 bl<60> cbl<30> in1<98> in2<98> sl<60> vdd vss wl<98> / cell_PIM
XI21944 bl<60> cbl<30> in1<97> in2<97> sl<60> vdd vss wl<97> / cell_PIM
XI21298 bl<52> cbl<26> in1<114> in2<114> sl<52> vdd vss wl<114> / cell_PIM
XI21297 bl<52> cbl<26> in1<113> in2<113> sl<52> vdd vss wl<113> / cell_PIM
XI21296 bl<52> cbl<26> in1<117> in2<117> sl<52> vdd vss wl<117> / cell_PIM
XI21295 bl<52> cbl<26> in1<116> in2<116> sl<52> vdd vss wl<116> / cell_PIM
XI22594 bl<36> cbl<18> in1<70> in2<70> sl<36> vdd vss wl<70> / cell_PIM
XI21289 bl<50> cbl<25> in1<113> in2<113> sl<50> vdd vss wl<113> / cell_PIM
XI21943 bl<60> cbl<30> in1<96> in2<96> sl<60> vdd vss wl<96> / cell_PIM
XI22592 bl<36> cbl<18> in1<73> in2<73> sl<36> vdd vss wl<73> / cell_PIM
XI22591 bl<36> cbl<18> in1<72> in2<72> sl<36> vdd vss wl<72> / cell_PIM
XI21288 bl<50> cbl<25> in1<114> in2<114> sl<50> vdd vss wl<114> / cell_PIM
XI21287 bl<50> cbl<25> in1<115> in2<115> sl<50> vdd vss wl<115> / cell_PIM
XI21286 bl<50> cbl<25> in1<117> in2<117> sl<50> vdd vss wl<117> / cell_PIM
XI21285 bl<50> cbl<25> in1<116> in2<116> sl<50> vdd vss wl<116> / cell_PIM
XI21937 bl<58> cbl<29> in1<94> in2<94> sl<58> vdd vss wl<94> / cell_PIM
XI21936 bl<58> cbl<29> in1<95> in2<95> sl<58> vdd vss wl<95> / cell_PIM
XI21935 bl<58> cbl<29> in1<97> in2<97> sl<58> vdd vss wl<97> / cell_PIM
XI21934 bl<58> cbl<29> in1<98> in2<98> sl<58> vdd vss wl<98> / cell_PIM
XI22585 bl<34> cbl<17> in1<70> in2<70> sl<34> vdd vss wl<70> / cell_PIM
XI22584 bl<34> cbl<17> in1<71> in2<71> sl<34> vdd vss wl<71> / cell_PIM
XI21279 bl<48> cbl<24> in1<115> in2<115> sl<48> vdd vss wl<115> / cell_PIM
XI21933 bl<58> cbl<29> in1<96> in2<96> sl<58> vdd vss wl<96> / cell_PIM
XI22582 bl<34> cbl<17> in1<74> in2<74> sl<34> vdd vss wl<74> / cell_PIM
XI22581 bl<34> cbl<17> in1<72> in2<72> sl<34> vdd vss wl<72> / cell_PIM
XI22575 bl<32> cbl<16> in1<71> in2<71> sl<32> vdd vss wl<71> / cell_PIM
XI21927 bl<56> cbl<28> in1<94> in2<94> sl<56> vdd vss wl<94> / cell_PIM
XI21926 bl<56> cbl<28> in1<95> in2<95> sl<56> vdd vss wl<95> / cell_PIM
XI21925 bl<56> cbl<28> in1<97> in2<97> sl<56> vdd vss wl<97> / cell_PIM
XI21924 bl<56> cbl<28> in1<98> in2<98> sl<56> vdd vss wl<98> / cell_PIM
XI21278 bl<48> cbl<24> in1<114> in2<114> sl<48> vdd vss wl<114> / cell_PIM
XI21277 bl<48> cbl<24> in1<113> in2<113> sl<48> vdd vss wl<113> / cell_PIM
XI21276 bl<48> cbl<24> in1<117> in2<117> sl<48> vdd vss wl<117> / cell_PIM
XI21275 bl<48> cbl<24> in1<116> in2<116> sl<48> vdd vss wl<116> / cell_PIM
XI22574 bl<32> cbl<16> in1<70> in2<70> sl<32> vdd vss wl<70> / cell_PIM
XI21269 bl<46> cbl<23> in1<113> in2<113> sl<46> vdd vss wl<113> / cell_PIM
XI21923 bl<56> cbl<28> in1<96> in2<96> sl<56> vdd vss wl<96> / cell_PIM
XI22572 bl<32> cbl<16> in1<73> in2<73> sl<32> vdd vss wl<73> / cell_PIM
XI22571 bl<32> cbl<16> in1<72> in2<72> sl<32> vdd vss wl<72> / cell_PIM
XI21268 bl<46> cbl<23> in1<114> in2<114> sl<46> vdd vss wl<114> / cell_PIM
XI21267 bl<46> cbl<23> in1<115> in2<115> sl<46> vdd vss wl<115> / cell_PIM
XI21266 bl<46> cbl<23> in1<117> in2<117> sl<46> vdd vss wl<117> / cell_PIM
XI21265 bl<46> cbl<23> in1<116> in2<116> sl<46> vdd vss wl<116> / cell_PIM
XI21917 bl<54> cbl<27> in1<94> in2<94> sl<54> vdd vss wl<94> / cell_PIM
XI21916 bl<54> cbl<27> in1<95> in2<95> sl<54> vdd vss wl<95> / cell_PIM
XI21915 bl<54> cbl<27> in1<97> in2<97> sl<54> vdd vss wl<97> / cell_PIM
XI21914 bl<54> cbl<27> in1<98> in2<98> sl<54> vdd vss wl<98> / cell_PIM
XI22565 bl<62> cbl<31> in1<75> in2<75> sl<62> vdd vss wl<75> / cell_PIM
XI22564 bl<62> cbl<31> in1<76> in2<76> sl<62> vdd vss wl<76> / cell_PIM
XI19759 bl<16> cbl<8> in1<67> in2<67> sl<16> vdd vss wl<67> / cell_PIM
XI20284 bl<16> cbl<8> in1<35> in2<35> sl<16> vdd vss wl<35> / cell_PIM
XI20283 bl<16> cbl<8> in1<34> in2<34> sl<16> vdd vss wl<34> / cell_PIM
XI20929 bl<42> cbl<21> in1<127> in2<127> sl<42> vdd vss wl<127> / cell_PIM
XI20928 bl<42> cbl<21> in1<126> in2<126> sl<42> vdd vss wl<126> / cell_PIM
XI20927 bl<42> cbl<21> in1<125> in2<125> sl<42> vdd vss wl<125> / cell_PIM
XI20926 bl<42> cbl<21> in1<123> in2<123> sl<42> vdd vss wl<123> / cell_PIM
XI20925 bl<42> cbl<21> in1<124> in2<124> sl<42> vdd vss wl<124> / cell_PIM
XI20278 bl<30> cbl<15> in1<37> in2<37> sl<30> vdd vss wl<37> / cell_PIM
XI20277 bl<30> cbl<15> in1<38> in2<38> sl<30> vdd vss wl<38> / cell_PIM
XI19758 bl<16> cbl<8> in1<66> in2<66> sl<16> vdd vss wl<66> / cell_PIM
XI19757 bl<16> cbl<8> in1<65> in2<65> sl<16> vdd vss wl<65> / cell_PIM
XI19756 bl<16> cbl<8> in1<69> in2<69> sl<16> vdd vss wl<69> / cell_PIM
XI19755 bl<16> cbl<8> in1<68> in2<68> sl<16> vdd vss wl<68> / cell_PIM
XI19749 bl<30> cbl<15> in1<70> in2<70> sl<30> vdd vss wl<70> / cell_PIM
XI20276 bl<30> cbl<15> in1<40> in2<40> sl<30> vdd vss wl<40> / cell_PIM
XI20275 bl<30> cbl<15> in1<39> in2<39> sl<30> vdd vss wl<39> / cell_PIM
XI20919 bl<40> cbl<20> in1<127> in2<127> sl<40> vdd vss wl<127> / cell_PIM
XI19747 bl<30> cbl<15> in1<73> in2<73> sl<30> vdd vss wl<73> / cell_PIM
XI19746 bl<30> cbl<15> in1<74> in2<74> sl<30> vdd vss wl<74> / cell_PIM
XI19745 bl<30> cbl<15> in1<72> in2<72> sl<30> vdd vss wl<72> / cell_PIM
XI19748 bl<30> cbl<15> in1<71> in2<71> sl<30> vdd vss wl<71> / cell_PIM
XI20270 bl<28> cbl<14> in1<38> in2<38> sl<28> vdd vss wl<38> / cell_PIM
XI20269 bl<28> cbl<14> in1<37> in2<37> sl<28> vdd vss wl<37> / cell_PIM
XI20918 bl<40> cbl<20> in1<126> in2<126> sl<40> vdd vss wl<126> / cell_PIM
XI20917 bl<40> cbl<20> in1<125> in2<125> sl<40> vdd vss wl<125> / cell_PIM
XI20916 bl<40> cbl<20> in1<123> in2<123> sl<40> vdd vss wl<123> / cell_PIM
XI20915 bl<40> cbl<20> in1<124> in2<124> sl<40> vdd vss wl<124> / cell_PIM
XI19739 bl<28> cbl<14> in1<71> in2<71> sl<28> vdd vss wl<71> / cell_PIM
XI20268 bl<28> cbl<14> in1<40> in2<40> sl<28> vdd vss wl<40> / cell_PIM
XI20267 bl<28> cbl<14> in1<39> in2<39> sl<28> vdd vss wl<39> / cell_PIM
XI20909 bl<38> cbl<19> in1<127> in2<127> sl<38> vdd vss wl<127> / cell_PIM
XI20908 bl<38> cbl<19> in1<126> in2<126> sl<38> vdd vss wl<126> / cell_PIM
XI20907 bl<38> cbl<19> in1<125> in2<125> sl<38> vdd vss wl<125> / cell_PIM
XI20906 bl<38> cbl<19> in1<123> in2<123> sl<38> vdd vss wl<123> / cell_PIM
XI20905 bl<38> cbl<19> in1<124> in2<124> sl<38> vdd vss wl<124> / cell_PIM
XI20262 bl<26> cbl<13> in1<37> in2<37> sl<26> vdd vss wl<37> / cell_PIM
XI20261 bl<26> cbl<13> in1<38> in2<38> sl<26> vdd vss wl<38> / cell_PIM
XI19738 bl<28> cbl<14> in1<70> in2<70> sl<28> vdd vss wl<70> / cell_PIM
XI19737 bl<28> cbl<14> in1<74> in2<74> sl<28> vdd vss wl<74> / cell_PIM
XI19736 bl<28> cbl<14> in1<73> in2<73> sl<28> vdd vss wl<73> / cell_PIM
XI19735 bl<28> cbl<14> in1<72> in2<72> sl<28> vdd vss wl<72> / cell_PIM
XI19729 bl<26> cbl<13> in1<70> in2<70> sl<26> vdd vss wl<70> / cell_PIM
XI20260 bl<26> cbl<13> in1<40> in2<40> sl<26> vdd vss wl<40> / cell_PIM
XI20259 bl<26> cbl<13> in1<39> in2<39> sl<26> vdd vss wl<39> / cell_PIM
XI20899 bl<36> cbl<18> in1<127> in2<127> sl<36> vdd vss wl<127> / cell_PIM
XI19727 bl<26> cbl<13> in1<73> in2<73> sl<26> vdd vss wl<73> / cell_PIM
XI19726 bl<26> cbl<13> in1<74> in2<74> sl<26> vdd vss wl<74> / cell_PIM
XI19725 bl<26> cbl<13> in1<72> in2<72> sl<26> vdd vss wl<72> / cell_PIM
XI19728 bl<26> cbl<13> in1<71> in2<71> sl<26> vdd vss wl<71> / cell_PIM
XI20254 bl<24> cbl<12> in1<37> in2<37> sl<24> vdd vss wl<37> / cell_PIM
XI20253 bl<24> cbl<12> in1<38> in2<38> sl<24> vdd vss wl<38> / cell_PIM
XI20898 bl<36> cbl<18> in1<126> in2<126> sl<36> vdd vss wl<126> / cell_PIM
XI20897 bl<36> cbl<18> in1<125> in2<125> sl<36> vdd vss wl<125> / cell_PIM
XI20896 bl<36> cbl<18> in1<124> in2<124> sl<36> vdd vss wl<124> / cell_PIM
XI20895 bl<36> cbl<18> in1<123> in2<123> sl<36> vdd vss wl<123> / cell_PIM
XI19719 bl<24> cbl<12> in1<70> in2<70> sl<24> vdd vss wl<70> / cell_PIM
XI20252 bl<24> cbl<12> in1<40> in2<40> sl<24> vdd vss wl<40> / cell_PIM
XI20251 bl<24> cbl<12> in1<39> in2<39> sl<24> vdd vss wl<39> / cell_PIM
XI20889 bl<34> cbl<17> in1<127> in2<127> sl<34> vdd vss wl<127> / cell_PIM
XI20888 bl<34> cbl<17> in1<126> in2<126> sl<34> vdd vss wl<126> / cell_PIM
XI20887 bl<34> cbl<17> in1<125> in2<125> sl<34> vdd vss wl<125> / cell_PIM
XI20886 bl<34> cbl<17> in1<123> in2<123> sl<34> vdd vss wl<123> / cell_PIM
XI20885 bl<34> cbl<17> in1<124> in2<124> sl<34> vdd vss wl<124> / cell_PIM
XI20246 bl<22> cbl<11> in1<37> in2<37> sl<22> vdd vss wl<37> / cell_PIM
XI20245 bl<22> cbl<11> in1<38> in2<38> sl<22> vdd vss wl<38> / cell_PIM
XI19718 bl<24> cbl<12> in1<71> in2<71> sl<24> vdd vss wl<71> / cell_PIM
XI19717 bl<24> cbl<12> in1<73> in2<73> sl<24> vdd vss wl<73> / cell_PIM
XI19716 bl<24> cbl<12> in1<74> in2<74> sl<24> vdd vss wl<74> / cell_PIM
XI19715 bl<24> cbl<12> in1<72> in2<72> sl<24> vdd vss wl<72> / cell_PIM
XI19709 bl<22> cbl<11> in1<70> in2<70> sl<22> vdd vss wl<70> / cell_PIM
XI20244 bl<22> cbl<11> in1<40> in2<40> sl<22> vdd vss wl<40> / cell_PIM
XI20243 bl<22> cbl<11> in1<39> in2<39> sl<22> vdd vss wl<39> / cell_PIM
XI20879 bl<32> cbl<16> in1<127> in2<127> sl<32> vdd vss wl<127> / cell_PIM
XI19707 bl<22> cbl<11> in1<73> in2<73> sl<22> vdd vss wl<73> / cell_PIM
XI19706 bl<22> cbl<11> in1<74> in2<74> sl<22> vdd vss wl<74> / cell_PIM
XI19705 bl<22> cbl<11> in1<72> in2<72> sl<22> vdd vss wl<72> / cell_PIM
XI19708 bl<22> cbl<11> in1<71> in2<71> sl<22> vdd vss wl<71> / cell_PIM
XI20238 bl<20> cbl<10> in1<38> in2<38> sl<20> vdd vss wl<38> / cell_PIM
XI20237 bl<20> cbl<10> in1<37> in2<37> sl<20> vdd vss wl<37> / cell_PIM
XI20878 bl<32> cbl<16> in1<126> in2<126> sl<32> vdd vss wl<126> / cell_PIM
XI20877 bl<32> cbl<16> in1<125> in2<125> sl<32> vdd vss wl<125> / cell_PIM
XI20876 bl<32> cbl<16> in1<124> in2<124> sl<32> vdd vss wl<124> / cell_PIM
XI20875 bl<32> cbl<16> in1<123> in2<123> sl<32> vdd vss wl<123> / cell_PIM
XI19699 bl<20> cbl<10> in1<71> in2<71> sl<20> vdd vss wl<71> / cell_PIM
XI20236 bl<20> cbl<10> in1<40> in2<40> sl<20> vdd vss wl<40> / cell_PIM
XI20235 bl<20> cbl<10> in1<39> in2<39> sl<20> vdd vss wl<39> / cell_PIM
XI20871 bl<30> cbl<15> in1<0> in2<0> sl<30> vdd vss wl<0> / cell_PIM
XI20870 bl<30> cbl<15> in1<1> in2<1> sl<30> vdd vss wl<1> / cell_PIM
XI20869 bl<30> cbl<15> in1<2> in2<2> sl<30> vdd vss wl<2> / cell_PIM
XI20865 bl<28> cbl<14> in1<0> in2<0> sl<28> vdd vss wl<0> / cell_PIM
XI20864 bl<28> cbl<14> in1<2> in2<2> sl<28> vdd vss wl<2> / cell_PIM
XI20230 bl<18> cbl<9> in1<37> in2<37> sl<18> vdd vss wl<37> / cell_PIM
XI20229 bl<18> cbl<9> in1<38> in2<38> sl<18> vdd vss wl<38> / cell_PIM
XI19698 bl<20> cbl<10> in1<70> in2<70> sl<20> vdd vss wl<70> / cell_PIM
XI19697 bl<20> cbl<10> in1<74> in2<74> sl<20> vdd vss wl<74> / cell_PIM
XI19696 bl<20> cbl<10> in1<73> in2<73> sl<20> vdd vss wl<73> / cell_PIM
XI19695 bl<20> cbl<10> in1<72> in2<72> sl<20> vdd vss wl<72> / cell_PIM
XI19689 bl<18> cbl<9> in1<70> in2<70> sl<18> vdd vss wl<70> / cell_PIM
XI20228 bl<18> cbl<9> in1<40> in2<40> sl<18> vdd vss wl<40> / cell_PIM
XI20227 bl<18> cbl<9> in1<39> in2<39> sl<18> vdd vss wl<39> / cell_PIM
XI20863 bl<28> cbl<14> in1<1> in2<1> sl<28> vdd vss wl<1> / cell_PIM
XI20859 bl<26> cbl<13> in1<0> in2<0> sl<26> vdd vss wl<0> / cell_PIM
XI19687 bl<18> cbl<9> in1<73> in2<73> sl<18> vdd vss wl<73> / cell_PIM
XI19686 bl<18> cbl<9> in1<74> in2<74> sl<18> vdd vss wl<74> / cell_PIM
XI19685 bl<18> cbl<9> in1<72> in2<72> sl<18> vdd vss wl<72> / cell_PIM
XI19688 bl<18> cbl<9> in1<71> in2<71> sl<18> vdd vss wl<71> / cell_PIM
XI20222 bl<16> cbl<8> in1<38> in2<38> sl<16> vdd vss wl<38> / cell_PIM
XI20221 bl<16> cbl<8> in1<37> in2<37> sl<16> vdd vss wl<37> / cell_PIM
XI20858 bl<26> cbl<13> in1<1> in2<1> sl<26> vdd vss wl<1> / cell_PIM
XI20857 bl<26> cbl<13> in1<2> in2<2> sl<26> vdd vss wl<2> / cell_PIM
XI19679 bl<16> cbl<8> in1<71> in2<71> sl<16> vdd vss wl<71> / cell_PIM
XI20220 bl<16> cbl<8> in1<40> in2<40> sl<16> vdd vss wl<40> / cell_PIM
XI20219 bl<16> cbl<8> in1<39> in2<39> sl<16> vdd vss wl<39> / cell_PIM
XI20853 bl<24> cbl<12> in1<0> in2<0> sl<24> vdd vss wl<0> / cell_PIM
XI20852 bl<24> cbl<12> in1<2> in2<2> sl<24> vdd vss wl<2> / cell_PIM
XI20851 bl<24> cbl<12> in1<1> in2<1> sl<24> vdd vss wl<1> / cell_PIM
XI20847 bl<22> cbl<11> in1<0> in2<0> sl<22> vdd vss wl<0> / cell_PIM
XI20846 bl<22> cbl<11> in1<1> in2<1> sl<22> vdd vss wl<1> / cell_PIM
XI20845 bl<22> cbl<11> in1<2> in2<2> sl<22> vdd vss wl<2> / cell_PIM
XI20213 bl<30> cbl<15> in1<41> in2<41> sl<30> vdd vss wl<41> / cell_PIM
XI19678 bl<16> cbl<8> in1<70> in2<70> sl<16> vdd vss wl<70> / cell_PIM
XI19677 bl<16> cbl<8> in1<74> in2<74> sl<16> vdd vss wl<74> / cell_PIM
XI19676 bl<16> cbl<8> in1<73> in2<73> sl<16> vdd vss wl<73> / cell_PIM
XI19675 bl<16> cbl<8> in1<72> in2<72> sl<16> vdd vss wl<72> / cell_PIM
XI19669 bl<30> cbl<15> in1<75> in2<75> sl<30> vdd vss wl<75> / cell_PIM
XI20212 bl<30> cbl<15> in1<42> in2<42> sl<30> vdd vss wl<42> / cell_PIM
XI20211 bl<30> cbl<15> in1<43> in2<43> sl<30> vdd vss wl<43> / cell_PIM
XI20210 bl<30> cbl<15> in1<45> in2<45> sl<30> vdd vss wl<45> / cell_PIM
XI20209 bl<30> cbl<15> in1<44> in2<44> sl<30> vdd vss wl<44> / cell_PIM
XI20841 bl<20> cbl<10> in1<0> in2<0> sl<20> vdd vss wl<0> / cell_PIM
XI20840 bl<20> cbl<10> in1<2> in2<2> sl<20> vdd vss wl<2> / cell_PIM
XI20839 bl<20> cbl<10> in1<1> in2<1> sl<20> vdd vss wl<1> / cell_PIM
XI19667 bl<30> cbl<15> in1<78> in2<78> sl<30> vdd vss wl<78> / cell_PIM
XI19666 bl<30> cbl<15> in1<79> in2<79> sl<30> vdd vss wl<79> / cell_PIM
XI19665 bl<30> cbl<15> in1<77> in2<77> sl<30> vdd vss wl<77> / cell_PIM
XI19668 bl<30> cbl<15> in1<76> in2<76> sl<30> vdd vss wl<76> / cell_PIM
XI20835 bl<18> cbl<9> in1<0> in2<0> sl<18> vdd vss wl<0> / cell_PIM
XI20834 bl<18> cbl<9> in1<1> in2<1> sl<18> vdd vss wl<1> / cell_PIM
XI19659 bl<28> cbl<14> in1<76> in2<76> sl<28> vdd vss wl<76> / cell_PIM
XI20203 bl<28> cbl<14> in1<43> in2<43> sl<28> vdd vss wl<43> / cell_PIM
XI20202 bl<28> cbl<14> in1<42> in2<42> sl<28> vdd vss wl<42> / cell_PIM
XI20201 bl<28> cbl<14> in1<41> in2<41> sl<28> vdd vss wl<41> / cell_PIM
XI20833 bl<18> cbl<9> in1<2> in2<2> sl<18> vdd vss wl<2> / cell_PIM
XI20829 bl<16> cbl<8> in1<0> in2<0> sl<16> vdd vss wl<0> / cell_PIM
XI20828 bl<16> cbl<8> in1<2> in2<2> sl<16> vdd vss wl<2> / cell_PIM
XI20827 bl<16> cbl<8> in1<1> in2<1> sl<16> vdd vss wl<1> / cell_PIM
XI20200 bl<28> cbl<14> in1<45> in2<45> sl<28> vdd vss wl<45> / cell_PIM
XI20199 bl<28> cbl<14> in1<44> in2<44> sl<28> vdd vss wl<44> / cell_PIM
XI19658 bl<28> cbl<14> in1<75> in2<75> sl<28> vdd vss wl<75> / cell_PIM
XI19657 bl<28> cbl<14> in1<79> in2<79> sl<28> vdd vss wl<79> / cell_PIM
XI19656 bl<28> cbl<14> in1<78> in2<78> sl<28> vdd vss wl<78> / cell_PIM
XI19655 bl<28> cbl<14> in1<77> in2<77> sl<28> vdd vss wl<77> / cell_PIM
XI19649 bl<26> cbl<13> in1<75> in2<75> sl<26> vdd vss wl<75> / cell_PIM
XI20193 bl<26> cbl<13> in1<41> in2<41> sl<26> vdd vss wl<41> / cell_PIM
XI20821 bl<30> cbl<15> in1<3> in2<3> sl<30> vdd vss wl<3> / cell_PIM
XI20820 bl<30> cbl<15> in1<4> in2<4> sl<30> vdd vss wl<4> / cell_PIM
XI20819 bl<30> cbl<15> in1<6> in2<6> sl<30> vdd vss wl<6> / cell_PIM
XI19647 bl<26> cbl<13> in1<78> in2<78> sl<26> vdd vss wl<78> / cell_PIM
XI19646 bl<26> cbl<13> in1<79> in2<79> sl<26> vdd vss wl<79> / cell_PIM
XI19645 bl<26> cbl<13> in1<77> in2<77> sl<26> vdd vss wl<77> / cell_PIM
XI19648 bl<26> cbl<13> in1<76> in2<76> sl<26> vdd vss wl<76> / cell_PIM
XI20192 bl<26> cbl<13> in1<42> in2<42> sl<26> vdd vss wl<42> / cell_PIM
XI20191 bl<26> cbl<13> in1<43> in2<43> sl<26> vdd vss wl<43> / cell_PIM
XI20190 bl<26> cbl<13> in1<45> in2<45> sl<26> vdd vss wl<45> / cell_PIM
XI20189 bl<26> cbl<13> in1<44> in2<44> sl<26> vdd vss wl<44> / cell_PIM
XI20818 bl<30> cbl<15> in1<7> in2<7> sl<30> vdd vss wl<7> / cell_PIM
XI20817 bl<30> cbl<15> in1<5> in2<5> sl<30> vdd vss wl<5> / cell_PIM
XI19639 bl<24> cbl<12> in1<75> in2<75> sl<24> vdd vss wl<75> / cell_PIM
XI20811 bl<28> cbl<14> in1<4> in2<4> sl<28> vdd vss wl<4> / cell_PIM
XI20810 bl<28> cbl<14> in1<3> in2<3> sl<28> vdd vss wl<3> / cell_PIM
XI20809 bl<28> cbl<14> in1<7> in2<7> sl<28> vdd vss wl<7> / cell_PIM
XI20808 bl<28> cbl<14> in1<6> in2<6> sl<28> vdd vss wl<6> / cell_PIM
XI20807 bl<28> cbl<14> in1<5> in2<5> sl<28> vdd vss wl<5> / cell_PIM
XI20183 bl<24> cbl<12> in1<41> in2<41> sl<24> vdd vss wl<41> / cell_PIM
XI20182 bl<24> cbl<12> in1<42> in2<42> sl<24> vdd vss wl<42> / cell_PIM
XI20181 bl<24> cbl<12> in1<43> in2<43> sl<24> vdd vss wl<43> / cell_PIM
XI19638 bl<24> cbl<12> in1<76> in2<76> sl<24> vdd vss wl<76> / cell_PIM
XI19637 bl<24> cbl<12> in1<78> in2<78> sl<24> vdd vss wl<78> / cell_PIM
XI19636 bl<24> cbl<12> in1<79> in2<79> sl<24> vdd vss wl<79> / cell_PIM
XI19635 bl<24> cbl<12> in1<77> in2<77> sl<24> vdd vss wl<77> / cell_PIM
XI19629 bl<22> cbl<11> in1<75> in2<75> sl<22> vdd vss wl<75> / cell_PIM
XI20180 bl<24> cbl<12> in1<45> in2<45> sl<24> vdd vss wl<45> / cell_PIM
XI20179 bl<24> cbl<12> in1<44> in2<44> sl<24> vdd vss wl<44> / cell_PIM
XI20801 bl<26> cbl<13> in1<3> in2<3> sl<26> vdd vss wl<3> / cell_PIM
XI20800 bl<26> cbl<13> in1<4> in2<4> sl<26> vdd vss wl<4> / cell_PIM
XI20799 bl<26> cbl<13> in1<6> in2<6> sl<26> vdd vss wl<6> / cell_PIM
XI19627 bl<22> cbl<11> in1<78> in2<78> sl<22> vdd vss wl<78> / cell_PIM
XI19626 bl<22> cbl<11> in1<79> in2<79> sl<22> vdd vss wl<79> / cell_PIM
XI19625 bl<22> cbl<11> in1<77> in2<77> sl<22> vdd vss wl<77> / cell_PIM
XI19628 bl<22> cbl<11> in1<76> in2<76> sl<22> vdd vss wl<76> / cell_PIM
XI20173 bl<22> cbl<11> in1<41> in2<41> sl<22> vdd vss wl<41> / cell_PIM
XI20798 bl<26> cbl<13> in1<7> in2<7> sl<26> vdd vss wl<7> / cell_PIM
XI20797 bl<26> cbl<13> in1<5> in2<5> sl<26> vdd vss wl<5> / cell_PIM
XI19619 bl<20> cbl<10> in1<76> in2<76> sl<20> vdd vss wl<76> / cell_PIM
XI20172 bl<22> cbl<11> in1<42> in2<42> sl<22> vdd vss wl<42> / cell_PIM
XI20171 bl<22> cbl<11> in1<43> in2<43> sl<22> vdd vss wl<43> / cell_PIM
XI20170 bl<22> cbl<11> in1<45> in2<45> sl<22> vdd vss wl<45> / cell_PIM
XI20169 bl<22> cbl<11> in1<44> in2<44> sl<22> vdd vss wl<44> / cell_PIM
XI20791 bl<24> cbl<12> in1<3> in2<3> sl<24> vdd vss wl<3> / cell_PIM
XI20790 bl<24> cbl<12> in1<4> in2<4> sl<24> vdd vss wl<4> / cell_PIM
XI20789 bl<24> cbl<12> in1<6> in2<6> sl<24> vdd vss wl<6> / cell_PIM
XI20788 bl<24> cbl<12> in1<7> in2<7> sl<24> vdd vss wl<7> / cell_PIM
XI20787 bl<24> cbl<12> in1<5> in2<5> sl<24> vdd vss wl<5> / cell_PIM
XI19618 bl<20> cbl<10> in1<75> in2<75> sl<20> vdd vss wl<75> / cell_PIM
XI19617 bl<20> cbl<10> in1<79> in2<79> sl<20> vdd vss wl<79> / cell_PIM
XI19616 bl<20> cbl<10> in1<78> in2<78> sl<20> vdd vss wl<78> / cell_PIM
XI19615 bl<20> cbl<10> in1<77> in2<77> sl<20> vdd vss wl<77> / cell_PIM
XI19609 bl<18> cbl<9> in1<75> in2<75> sl<18> vdd vss wl<75> / cell_PIM
XI20163 bl<20> cbl<10> in1<43> in2<43> sl<20> vdd vss wl<43> / cell_PIM
XI20162 bl<20> cbl<10> in1<42> in2<42> sl<20> vdd vss wl<42> / cell_PIM
XI20161 bl<20> cbl<10> in1<41> in2<41> sl<20> vdd vss wl<41> / cell_PIM
XI20781 bl<22> cbl<11> in1<3> in2<3> sl<22> vdd vss wl<3> / cell_PIM
XI20780 bl<22> cbl<11> in1<4> in2<4> sl<22> vdd vss wl<4> / cell_PIM
XI20779 bl<22> cbl<11> in1<6> in2<6> sl<22> vdd vss wl<6> / cell_PIM
XI19607 bl<18> cbl<9> in1<78> in2<78> sl<18> vdd vss wl<78> / cell_PIM
XI19606 bl<18> cbl<9> in1<79> in2<79> sl<18> vdd vss wl<79> / cell_PIM
XI19605 bl<18> cbl<9> in1<77> in2<77> sl<18> vdd vss wl<77> / cell_PIM
XI19608 bl<18> cbl<9> in1<76> in2<76> sl<18> vdd vss wl<76> / cell_PIM
XI20160 bl<20> cbl<10> in1<45> in2<45> sl<20> vdd vss wl<45> / cell_PIM
XI20159 bl<20> cbl<10> in1<44> in2<44> sl<20> vdd vss wl<44> / cell_PIM
XI20778 bl<22> cbl<11> in1<7> in2<7> sl<22> vdd vss wl<7> / cell_PIM
XI20777 bl<22> cbl<11> in1<5> in2<5> sl<22> vdd vss wl<5> / cell_PIM
XI19599 bl<16> cbl<8> in1<76> in2<76> sl<16> vdd vss wl<76> / cell_PIM
XI20153 bl<18> cbl<9> in1<41> in2<41> sl<18> vdd vss wl<41> / cell_PIM
XI20771 bl<20> cbl<10> in1<4> in2<4> sl<20> vdd vss wl<4> / cell_PIM
XI20770 bl<20> cbl<10> in1<3> in2<3> sl<20> vdd vss wl<3> / cell_PIM
XI20769 bl<20> cbl<10> in1<7> in2<7> sl<20> vdd vss wl<7> / cell_PIM
XI20768 bl<20> cbl<10> in1<6> in2<6> sl<20> vdd vss wl<6> / cell_PIM
XI20767 bl<20> cbl<10> in1<5> in2<5> sl<20> vdd vss wl<5> / cell_PIM
XI20152 bl<18> cbl<9> in1<42> in2<42> sl<18> vdd vss wl<42> / cell_PIM
XI20151 bl<18> cbl<9> in1<43> in2<43> sl<18> vdd vss wl<43> / cell_PIM
XI20150 bl<18> cbl<9> in1<45> in2<45> sl<18> vdd vss wl<45> / cell_PIM
XI20149 bl<18> cbl<9> in1<44> in2<44> sl<18> vdd vss wl<44> / cell_PIM
XI19598 bl<16> cbl<8> in1<75> in2<75> sl<16> vdd vss wl<75> / cell_PIM
XI19597 bl<16> cbl<8> in1<79> in2<79> sl<16> vdd vss wl<79> / cell_PIM
XI19596 bl<16> cbl<8> in1<78> in2<78> sl<16> vdd vss wl<78> / cell_PIM
XI19595 bl<16> cbl<8> in1<77> in2<77> sl<16> vdd vss wl<77> / cell_PIM
XI19590 bl<30> cbl<15> in1<80> in2<80> sl<30> vdd vss wl<80> / cell_PIM
XI19589 bl<30> cbl<15> in1<81> in2<81> sl<30> vdd vss wl<81> / cell_PIM
XI20761 bl<18> cbl<9> in1<3> in2<3> sl<18> vdd vss wl<3> / cell_PIM
XI20760 bl<18> cbl<9> in1<4> in2<4> sl<18> vdd vss wl<4> / cell_PIM
XI20759 bl<18> cbl<9> in1<6> in2<6> sl<18> vdd vss wl<6> / cell_PIM
XI19587 bl<30> cbl<15> in1<82> in2<82> sl<30> vdd vss wl<82> / cell_PIM
XI19588 bl<30> cbl<15> in1<83> in2<83> sl<30> vdd vss wl<83> / cell_PIM
XI20143 bl<16> cbl<8> in1<43> in2<43> sl<16> vdd vss wl<43> / cell_PIM
XI20142 bl<16> cbl<8> in1<42> in2<42> sl<16> vdd vss wl<42> / cell_PIM
XI20141 bl<16> cbl<8> in1<41> in2<41> sl<16> vdd vss wl<41> / cell_PIM
XI20758 bl<18> cbl<9> in1<7> in2<7> sl<18> vdd vss wl<7> / cell_PIM
XI20757 bl<18> cbl<9> in1<5> in2<5> sl<18> vdd vss wl<5> / cell_PIM
XI19582 bl<28> cbl<14> in1<81> in2<81> sl<28> vdd vss wl<81> / cell_PIM
XI19581 bl<28> cbl<14> in1<80> in2<80> sl<28> vdd vss wl<80> / cell_PIM
XI19580 bl<28> cbl<14> in1<83> in2<83> sl<28> vdd vss wl<83> / cell_PIM
XI19579 bl<28> cbl<14> in1<82> in2<82> sl<28> vdd vss wl<82> / cell_PIM
XI20140 bl<16> cbl<8> in1<45> in2<45> sl<16> vdd vss wl<45> / cell_PIM
XI20139 bl<16> cbl<8> in1<44> in2<44> sl<16> vdd vss wl<44> / cell_PIM
XI20751 bl<16> cbl<8> in1<4> in2<4> sl<16> vdd vss wl<4> / cell_PIM
XI20750 bl<16> cbl<8> in1<3> in2<3> sl<16> vdd vss wl<3> / cell_PIM
XI20749 bl<16> cbl<8> in1<7> in2<7> sl<16> vdd vss wl<7> / cell_PIM
XI20748 bl<16> cbl<8> in1<6> in2<6> sl<16> vdd vss wl<6> / cell_PIM
XI20747 bl<16> cbl<8> in1<5> in2<5> sl<16> vdd vss wl<5> / cell_PIM
XI20133 bl<30> cbl<15> in1<46> in2<46> sl<30> vdd vss wl<46> / cell_PIM
XI19574 bl<26> cbl<13> in1<80> in2<80> sl<26> vdd vss wl<80> / cell_PIM
XI19572 bl<26> cbl<13> in1<83> in2<83> sl<26> vdd vss wl<83> / cell_PIM
XI19571 bl<26> cbl<13> in1<82> in2<82> sl<26> vdd vss wl<82> / cell_PIM
XI19573 bl<26> cbl<13> in1<81> in2<81> sl<26> vdd vss wl<81> / cell_PIM
XI20132 bl<30> cbl<15> in1<47> in2<47> sl<30> vdd vss wl<47> / cell_PIM
XI20131 bl<30> cbl<15> in1<49> in2<49> sl<30> vdd vss wl<49> / cell_PIM
XI20130 bl<30> cbl<15> in1<50> in2<50> sl<30> vdd vss wl<50> / cell_PIM
XI20129 bl<30> cbl<15> in1<48> in2<48> sl<30> vdd vss wl<48> / cell_PIM
XI20741 bl<30> cbl<15> in1<8> in2<8> sl<30> vdd vss wl<8> / cell_PIM
XI20740 bl<30> cbl<15> in1<9> in2<9> sl<30> vdd vss wl<9> / cell_PIM
XI20739 bl<30> cbl<15> in1<11> in2<11> sl<30> vdd vss wl<11> / cell_PIM
XI19566 bl<24> cbl<12> in1<80> in2<80> sl<24> vdd vss wl<80> / cell_PIM
XI19565 bl<24> cbl<12> in1<81> in2<81> sl<24> vdd vss wl<81> / cell_PIM
XI19564 bl<24> cbl<12> in1<83> in2<83> sl<24> vdd vss wl<83> / cell_PIM
XI20738 bl<30> cbl<15> in1<12> in2<12> sl<30> vdd vss wl<12> / cell_PIM
XI20737 bl<30> cbl<15> in1<10> in2<10> sl<30> vdd vss wl<10> / cell_PIM
XI19563 bl<24> cbl<12> in1<82> in2<82> sl<24> vdd vss wl<82> / cell_PIM
XI20123 bl<28> cbl<14> in1<47> in2<47> sl<28> vdd vss wl<47> / cell_PIM
XI20122 bl<28> cbl<14> in1<46> in2<46> sl<28> vdd vss wl<46> / cell_PIM
XI20121 bl<28> cbl<14> in1<50> in2<50> sl<28> vdd vss wl<50> / cell_PIM
XI20731 bl<28> cbl<14> in1<9> in2<9> sl<28> vdd vss wl<9> / cell_PIM
XI20730 bl<28> cbl<14> in1<8> in2<8> sl<28> vdd vss wl<8> / cell_PIM
XI20729 bl<28> cbl<14> in1<12> in2<12> sl<28> vdd vss wl<12> / cell_PIM
XI20728 bl<28> cbl<14> in1<11> in2<11> sl<28> vdd vss wl<11> / cell_PIM
XI20727 bl<28> cbl<14> in1<10> in2<10> sl<28> vdd vss wl<10> / cell_PIM
XI20120 bl<28> cbl<14> in1<49> in2<49> sl<28> vdd vss wl<49> / cell_PIM
XI20119 bl<28> cbl<14> in1<48> in2<48> sl<28> vdd vss wl<48> / cell_PIM
XI19558 bl<22> cbl<11> in1<80> in2<80> sl<22> vdd vss wl<80> / cell_PIM
XI19557 bl<22> cbl<11> in1<81> in2<81> sl<22> vdd vss wl<81> / cell_PIM
XI19556 bl<22> cbl<11> in1<83> in2<83> sl<22> vdd vss wl<83> / cell_PIM
XI19555 bl<22> cbl<11> in1<82> in2<82> sl<22> vdd vss wl<82> / cell_PIM
XI19550 bl<20> cbl<10> in1<81> in2<81> sl<20> vdd vss wl<81> / cell_PIM
XI19549 bl<20> cbl<10> in1<80> in2<80> sl<20> vdd vss wl<80> / cell_PIM
XI20113 bl<26> cbl<13> in1<46> in2<46> sl<26> vdd vss wl<46> / cell_PIM
XI20721 bl<26> cbl<13> in1<8> in2<8> sl<26> vdd vss wl<8> / cell_PIM
XI20720 bl<26> cbl<13> in1<9> in2<9> sl<26> vdd vss wl<9> / cell_PIM
XI20719 bl<26> cbl<13> in1<11> in2<11> sl<26> vdd vss wl<11> / cell_PIM
XI19547 bl<20> cbl<10> in1<82> in2<82> sl<20> vdd vss wl<82> / cell_PIM
XI19548 bl<20> cbl<10> in1<83> in2<83> sl<20> vdd vss wl<83> / cell_PIM
XI20112 bl<26> cbl<13> in1<47> in2<47> sl<26> vdd vss wl<47> / cell_PIM
XI20111 bl<26> cbl<13> in1<49> in2<49> sl<26> vdd vss wl<49> / cell_PIM
XI20110 bl<26> cbl<13> in1<50> in2<50> sl<26> vdd vss wl<50> / cell_PIM
XI20109 bl<26> cbl<13> in1<48> in2<48> sl<26> vdd vss wl<48> / cell_PIM
XI20718 bl<26> cbl<13> in1<12> in2<12> sl<26> vdd vss wl<12> / cell_PIM
XI20717 bl<26> cbl<13> in1<10> in2<10> sl<26> vdd vss wl<10> / cell_PIM
XI19542 bl<18> cbl<9> in1<80> in2<80> sl<18> vdd vss wl<80> / cell_PIM
XI19541 bl<18> cbl<9> in1<81> in2<81> sl<18> vdd vss wl<81> / cell_PIM
XI19540 bl<18> cbl<9> in1<83> in2<83> sl<18> vdd vss wl<83> / cell_PIM
XI19539 bl<18> cbl<9> in1<82> in2<82> sl<18> vdd vss wl<82> / cell_PIM
XI20711 bl<24> cbl<12> in1<8> in2<8> sl<24> vdd vss wl<8> / cell_PIM
XI20710 bl<24> cbl<12> in1<9> in2<9> sl<24> vdd vss wl<9> / cell_PIM
XI20709 bl<24> cbl<12> in1<11> in2<11> sl<24> vdd vss wl<11> / cell_PIM
XI20708 bl<24> cbl<12> in1<12> in2<12> sl<24> vdd vss wl<12> / cell_PIM
XI20707 bl<24> cbl<12> in1<10> in2<10> sl<24> vdd vss wl<10> / cell_PIM
XI20103 bl<24> cbl<12> in1<46> in2<46> sl<24> vdd vss wl<46> / cell_PIM
XI20102 bl<24> cbl<12> in1<47> in2<47> sl<24> vdd vss wl<47> / cell_PIM
XI20101 bl<24> cbl<12> in1<49> in2<49> sl<24> vdd vss wl<49> / cell_PIM
XI19534 bl<16> cbl<8> in1<81> in2<81> sl<16> vdd vss wl<81> / cell_PIM
XI19532 bl<16> cbl<8> in1<83> in2<83> sl<16> vdd vss wl<83> / cell_PIM
XI19531 bl<16> cbl<8> in1<82> in2<82> sl<16> vdd vss wl<82> / cell_PIM
XI19533 bl<16> cbl<8> in1<80> in2<80> sl<16> vdd vss wl<80> / cell_PIM
XI20100 bl<24> cbl<12> in1<50> in2<50> sl<24> vdd vss wl<50> / cell_PIM
XI20099 bl<24> cbl<12> in1<48> in2<48> sl<24> vdd vss wl<48> / cell_PIM
XI20701 bl<22> cbl<11> in1<8> in2<8> sl<22> vdd vss wl<8> / cell_PIM
XI20700 bl<22> cbl<11> in1<9> in2<9> sl<22> vdd vss wl<9> / cell_PIM
XI20699 bl<22> cbl<11> in1<11> in2<11> sl<22> vdd vss wl<11> / cell_PIM
XI19525 bl<30> cbl<15> in1<84> in2<84> sl<30> vdd vss wl<84> / cell_PIM
XI19524 bl<30> cbl<15> in1<85> in2<85> sl<30> vdd vss wl<85> / cell_PIM
XI20093 bl<22> cbl<11> in1<46> in2<46> sl<22> vdd vss wl<46> / cell_PIM
XI20698 bl<22> cbl<11> in1<12> in2<12> sl<22> vdd vss wl<12> / cell_PIM
XI20697 bl<22> cbl<11> in1<10> in2<10> sl<22> vdd vss wl<10> / cell_PIM
XI19522 bl<30> cbl<15> in1<88> in2<88> sl<30> vdd vss wl<88> / cell_PIM
XI19521 bl<30> cbl<15> in1<87> in2<87> sl<30> vdd vss wl<87> / cell_PIM
XI19523 bl<30> cbl<15> in1<86> in2<86> sl<30> vdd vss wl<86> / cell_PIM
XI20092 bl<22> cbl<11> in1<47> in2<47> sl<22> vdd vss wl<47> / cell_PIM
XI20091 bl<22> cbl<11> in1<49> in2<49> sl<22> vdd vss wl<49> / cell_PIM
XI20090 bl<22> cbl<11> in1<50> in2<50> sl<22> vdd vss wl<50> / cell_PIM
XI20089 bl<22> cbl<11> in1<48> in2<48> sl<22> vdd vss wl<48> / cell_PIM
XI20691 bl<20> cbl<10> in1<9> in2<9> sl<20> vdd vss wl<9> / cell_PIM
XI20690 bl<20> cbl<10> in1<8> in2<8> sl<20> vdd vss wl<8> / cell_PIM
XI20689 bl<20> cbl<10> in1<12> in2<12> sl<20> vdd vss wl<12> / cell_PIM
XI20688 bl<20> cbl<10> in1<11> in2<11> sl<20> vdd vss wl<11> / cell_PIM
XI20687 bl<20> cbl<10> in1<10> in2<10> sl<20> vdd vss wl<10> / cell_PIM
XI19515 bl<28> cbl<14> in1<86> in2<86> sl<28> vdd vss wl<86> / cell_PIM
XI19514 bl<28> cbl<14> in1<85> in2<85> sl<28> vdd vss wl<85> / cell_PIM
XI19512 bl<28> cbl<14> in1<88> in2<88> sl<28> vdd vss wl<88> / cell_PIM
XI19511 bl<28> cbl<14> in1<87> in2<87> sl<28> vdd vss wl<87> / cell_PIM
XI19513 bl<28> cbl<14> in1<84> in2<84> sl<28> vdd vss wl<84> / cell_PIM
XI20083 bl<20> cbl<10> in1<47> in2<47> sl<20> vdd vss wl<47> / cell_PIM
XI20082 bl<20> cbl<10> in1<46> in2<46> sl<20> vdd vss wl<46> / cell_PIM
XI20081 bl<20> cbl<10> in1<50> in2<50> sl<20> vdd vss wl<50> / cell_PIM
XI20681 bl<18> cbl<9> in1<8> in2<8> sl<18> vdd vss wl<8> / cell_PIM
XI20680 bl<18> cbl<9> in1<9> in2<9> sl<18> vdd vss wl<9> / cell_PIM
XI20679 bl<18> cbl<9> in1<11> in2<11> sl<18> vdd vss wl<11> / cell_PIM
XI19505 bl<26> cbl<13> in1<84> in2<84> sl<26> vdd vss wl<84> / cell_PIM
XI19504 bl<26> cbl<13> in1<85> in2<85> sl<26> vdd vss wl<85> / cell_PIM
XI20080 bl<20> cbl<10> in1<49> in2<49> sl<20> vdd vss wl<49> / cell_PIM
XI20079 bl<20> cbl<10> in1<48> in2<48> sl<20> vdd vss wl<48> / cell_PIM
XI20678 bl<18> cbl<9> in1<12> in2<12> sl<18> vdd vss wl<12> / cell_PIM
XI20677 bl<18> cbl<9> in1<10> in2<10> sl<18> vdd vss wl<10> / cell_PIM
XI19502 bl<26> cbl<13> in1<88> in2<88> sl<26> vdd vss wl<88> / cell_PIM
XI19501 bl<26> cbl<13> in1<87> in2<87> sl<26> vdd vss wl<87> / cell_PIM
XI19503 bl<26> cbl<13> in1<86> in2<86> sl<26> vdd vss wl<86> / cell_PIM
XI20073 bl<18> cbl<9> in1<46> in2<46> sl<18> vdd vss wl<46> / cell_PIM
XI20671 bl<16> cbl<8> in1<9> in2<9> sl<16> vdd vss wl<9> / cell_PIM
XI20670 bl<16> cbl<8> in1<8> in2<8> sl<16> vdd vss wl<8> / cell_PIM
XI20669 bl<16> cbl<8> in1<12> in2<12> sl<16> vdd vss wl<12> / cell_PIM
XI20668 bl<16> cbl<8> in1<11> in2<11> sl<16> vdd vss wl<11> / cell_PIM
XI20667 bl<16> cbl<8> in1<10> in2<10> sl<16> vdd vss wl<10> / cell_PIM
XI20072 bl<18> cbl<9> in1<47> in2<47> sl<18> vdd vss wl<47> / cell_PIM
XI20071 bl<18> cbl<9> in1<49> in2<49> sl<18> vdd vss wl<49> / cell_PIM
XI20070 bl<18> cbl<9> in1<50> in2<50> sl<18> vdd vss wl<50> / cell_PIM
XI20069 bl<18> cbl<9> in1<48> in2<48> sl<18> vdd vss wl<48> / cell_PIM
XI19495 bl<24> cbl<12> in1<84> in2<84> sl<24> vdd vss wl<84> / cell_PIM
XI19494 bl<24> cbl<12> in1<85> in2<85> sl<24> vdd vss wl<85> / cell_PIM
XI19492 bl<24> cbl<12> in1<88> in2<88> sl<24> vdd vss wl<88> / cell_PIM
XI19491 bl<24> cbl<12> in1<87> in2<87> sl<24> vdd vss wl<87> / cell_PIM
XI19493 bl<24> cbl<12> in1<86> in2<86> sl<24> vdd vss wl<86> / cell_PIM
XI20661 bl<30> cbl<15> in1<13> in2<13> sl<30> vdd vss wl<13> / cell_PIM
XI20660 bl<30> cbl<15> in1<14> in2<14> sl<30> vdd vss wl<14> / cell_PIM
XI20659 bl<30> cbl<15> in1<16> in2<16> sl<30> vdd vss wl<16> / cell_PIM
XI19485 bl<22> cbl<11> in1<84> in2<84> sl<22> vdd vss wl<84> / cell_PIM
XI19484 bl<22> cbl<11> in1<85> in2<85> sl<22> vdd vss wl<85> / cell_PIM
XI20063 bl<16> cbl<8> in1<47> in2<47> sl<16> vdd vss wl<47> / cell_PIM
XI20062 bl<16> cbl<8> in1<46> in2<46> sl<16> vdd vss wl<46> / cell_PIM
XI20061 bl<16> cbl<8> in1<50> in2<50> sl<16> vdd vss wl<50> / cell_PIM
XI20658 bl<30> cbl<15> in1<17> in2<17> sl<30> vdd vss wl<17> / cell_PIM
XI20657 bl<30> cbl<15> in1<15> in2<15> sl<30> vdd vss wl<15> / cell_PIM
XI19482 bl<22> cbl<11> in1<88> in2<88> sl<22> vdd vss wl<88> / cell_PIM
XI19481 bl<22> cbl<11> in1<87> in2<87> sl<22> vdd vss wl<87> / cell_PIM
XI19483 bl<22> cbl<11> in1<86> in2<86> sl<22> vdd vss wl<86> / cell_PIM
XI20060 bl<16> cbl<8> in1<49> in2<49> sl<16> vdd vss wl<49> / cell_PIM
XI20059 bl<16> cbl<8> in1<48> in2<48> sl<16> vdd vss wl<48> / cell_PIM
XI20651 bl<28> cbl<14> in1<14> in2<14> sl<28> vdd vss wl<14> / cell_PIM
XI20650 bl<28> cbl<14> in1<13> in2<13> sl<28> vdd vss wl<13> / cell_PIM
XI20649 bl<28> cbl<14> in1<17> in2<17> sl<28> vdd vss wl<17> / cell_PIM
XI20648 bl<28> cbl<14> in1<16> in2<16> sl<28> vdd vss wl<16> / cell_PIM
XI20647 bl<28> cbl<14> in1<15> in2<15> sl<28> vdd vss wl<15> / cell_PIM
XI20053 bl<30> cbl<15> in1<51> in2<51> sl<30> vdd vss wl<51> / cell_PIM
XI19475 bl<20> cbl<10> in1<86> in2<86> sl<20> vdd vss wl<86> / cell_PIM
XI19474 bl<20> cbl<10> in1<85> in2<85> sl<20> vdd vss wl<85> / cell_PIM
XI19472 bl<20> cbl<10> in1<88> in2<88> sl<20> vdd vss wl<88> / cell_PIM
XI19471 bl<20> cbl<10> in1<87> in2<87> sl<20> vdd vss wl<87> / cell_PIM
XI19473 bl<20> cbl<10> in1<84> in2<84> sl<20> vdd vss wl<84> / cell_PIM
XI20052 bl<30> cbl<15> in1<52> in2<52> sl<30> vdd vss wl<52> / cell_PIM
XI20051 bl<30> cbl<15> in1<54> in2<54> sl<30> vdd vss wl<54> / cell_PIM
XI20050 bl<30> cbl<15> in1<55> in2<55> sl<30> vdd vss wl<55> / cell_PIM
XI20049 bl<30> cbl<15> in1<53> in2<53> sl<30> vdd vss wl<53> / cell_PIM
XI20641 bl<26> cbl<13> in1<13> in2<13> sl<26> vdd vss wl<13> / cell_PIM
XI20640 bl<26> cbl<13> in1<14> in2<14> sl<26> vdd vss wl<14> / cell_PIM
XI20639 bl<26> cbl<13> in1<16> in2<16> sl<26> vdd vss wl<16> / cell_PIM
XI19465 bl<18> cbl<9> in1<84> in2<84> sl<18> vdd vss wl<84> / cell_PIM
XI19464 bl<18> cbl<9> in1<85> in2<85> sl<18> vdd vss wl<85> / cell_PIM
XI20638 bl<26> cbl<13> in1<17> in2<17> sl<26> vdd vss wl<17> / cell_PIM
XI20637 bl<26> cbl<13> in1<15> in2<15> sl<26> vdd vss wl<15> / cell_PIM
XI19462 bl<18> cbl<9> in1<88> in2<88> sl<18> vdd vss wl<88> / cell_PIM
XI19461 bl<18> cbl<9> in1<87> in2<87> sl<18> vdd vss wl<87> / cell_PIM
XI19463 bl<18> cbl<9> in1<86> in2<86> sl<18> vdd vss wl<86> / cell_PIM
XI20043 bl<28> cbl<14> in1<52> in2<52> sl<28> vdd vss wl<52> / cell_PIM
XI20042 bl<28> cbl<14> in1<51> in2<51> sl<28> vdd vss wl<51> / cell_PIM
XI20041 bl<28> cbl<14> in1<55> in2<55> sl<28> vdd vss wl<55> / cell_PIM
XI20631 bl<24> cbl<12> in1<13> in2<13> sl<24> vdd vss wl<13> / cell_PIM
XI20630 bl<24> cbl<12> in1<14> in2<14> sl<24> vdd vss wl<14> / cell_PIM
XI20629 bl<24> cbl<12> in1<16> in2<16> sl<24> vdd vss wl<16> / cell_PIM
XI20628 bl<24> cbl<12> in1<17> in2<17> sl<24> vdd vss wl<17> / cell_PIM
XI20627 bl<24> cbl<12> in1<15> in2<15> sl<24> vdd vss wl<15> / cell_PIM
XI20040 bl<28> cbl<14> in1<54> in2<54> sl<28> vdd vss wl<54> / cell_PIM
XI20039 bl<28> cbl<14> in1<53> in2<53> sl<28> vdd vss wl<53> / cell_PIM
XI19455 bl<16> cbl<8> in1<86> in2<86> sl<16> vdd vss wl<86> / cell_PIM
XI19454 bl<16> cbl<8> in1<85> in2<85> sl<16> vdd vss wl<85> / cell_PIM
XI19452 bl<16> cbl<8> in1<88> in2<88> sl<16> vdd vss wl<88> / cell_PIM
XI19451 bl<16> cbl<8> in1<87> in2<87> sl<16> vdd vss wl<87> / cell_PIM
XI19453 bl<16> cbl<8> in1<84> in2<84> sl<16> vdd vss wl<84> / cell_PIM
XI20033 bl<26> cbl<13> in1<51> in2<51> sl<26> vdd vss wl<51> / cell_PIM
XI20621 bl<22> cbl<11> in1<13> in2<13> sl<22> vdd vss wl<13> / cell_PIM
XI20620 bl<22> cbl<11> in1<14> in2<14> sl<22> vdd vss wl<14> / cell_PIM
XI20619 bl<22> cbl<11> in1<16> in2<16> sl<22> vdd vss wl<16> / cell_PIM
XI19445 bl<30> cbl<15> in1<89> in2<89> sl<30> vdd vss wl<89> / cell_PIM
XI19444 bl<30> cbl<15> in1<90> in2<90> sl<30> vdd vss wl<90> / cell_PIM
XI20032 bl<26> cbl<13> in1<52> in2<52> sl<26> vdd vss wl<52> / cell_PIM
XI20031 bl<26> cbl<13> in1<54> in2<54> sl<26> vdd vss wl<54> / cell_PIM
XI20030 bl<26> cbl<13> in1<55> in2<55> sl<26> vdd vss wl<55> / cell_PIM
XI20029 bl<26> cbl<13> in1<53> in2<53> sl<26> vdd vss wl<53> / cell_PIM
XI20618 bl<22> cbl<11> in1<17> in2<17> sl<22> vdd vss wl<17> / cell_PIM
XI20617 bl<22> cbl<11> in1<15> in2<15> sl<22> vdd vss wl<15> / cell_PIM
XI17811 bl<10> cbl<5> in1<127> in2<127> sl<10> vdd vss wl<127> / cell_PIM
XI17810 bl<10> cbl<5> in1<126> in2<126> sl<10> vdd vss wl<126> / cell_PIM
XI17809 bl<10> cbl<5> in1<125> in2<125> sl<10> vdd vss wl<125> / cell_PIM
XI18462 bl<12> cbl<6> in1<47> in2<47> sl<12> vdd vss wl<47> / cell_PIM
XI18461 bl<12> cbl<6> in1<46> in2<46> sl<12> vdd vss wl<46> / cell_PIM
XI18460 bl<12> cbl<6> in1<45> in2<45> sl<12> vdd vss wl<45> / cell_PIM
XI18459 bl<12> cbl<6> in1<44> in2<44> sl<12> vdd vss wl<44> / cell_PIM
XI19111 bl<24> cbl<12> in1<108> in2<108> sl<24> vdd vss wl<108> / cell_PIM
XI19110 bl<24> cbl<12> in1<109> in2<109> sl<24> vdd vss wl<109> / cell_PIM
XI19109 bl<24> cbl<12> in1<110> in2<110> sl<24> vdd vss wl<110> / cell_PIM
XI19108 bl<24> cbl<12> in1<112> in2<112> sl<24> vdd vss wl<112> / cell_PIM
XI19107 bl<24> cbl<12> in1<111> in2<111> sl<24> vdd vss wl<111> / cell_PIM
XI18454 bl<10> cbl<5> in1<45> in2<45> sl<10> vdd vss wl<45> / cell_PIM
XI17805 bl<8> cbl<4> in1<127> in2<127> sl<8> vdd vss wl<127> / cell_PIM
XI17804 bl<8> cbl<4> in1<126> in2<126> sl<8> vdd vss wl<126> / cell_PIM
XI17803 bl<8> cbl<4> in1<125> in2<125> sl<8> vdd vss wl<125> / cell_PIM
XI17801 bl<6> cbl<3> in1<0> in2<0> sl<6> vdd vss wl<0> / cell_PIM
XI17799 bl<4> cbl<2> in1<0> in2<0> sl<4> vdd vss wl<0> / cell_PIM
XI18453 bl<10> cbl<5> in1<46> in2<46> sl<10> vdd vss wl<46> / cell_PIM
XI18452 bl<10> cbl<5> in1<47> in2<47> sl<10> vdd vss wl<47> / cell_PIM
XI18451 bl<10> cbl<5> in1<44> in2<44> sl<10> vdd vss wl<44> / cell_PIM
XI19101 bl<22> cbl<11> in1<108> in2<108> sl<22> vdd vss wl<108> / cell_PIM
XI19100 bl<22> cbl<11> in1<109> in2<109> sl<22> vdd vss wl<109> / cell_PIM
XI19099 bl<22> cbl<11> in1<110> in2<110> sl<22> vdd vss wl<110> / cell_PIM
XI17794 bl<6> cbl<3> in1<1> in2<1> sl<6> vdd vss wl<1> / cell_PIM
XI18446 bl<8> cbl<4> in1<47> in2<47> sl<8> vdd vss wl<47> / cell_PIM
XI18445 bl<8> cbl<4> in1<46> in2<46> sl<8> vdd vss wl<46> / cell_PIM
XI18444 bl<8> cbl<4> in1<45> in2<45> sl<8> vdd vss wl<45> / cell_PIM
XI19098 bl<22> cbl<11> in1<112> in2<112> sl<22> vdd vss wl<112> / cell_PIM
XI19097 bl<22> cbl<11> in1<111> in2<111> sl<22> vdd vss wl<111> / cell_PIM
XI17793 bl<6> cbl<3> in1<2> in2<2> sl<6> vdd vss wl<2> / cell_PIM
XI17792 bl<6> cbl<3> in1<3> in2<3> sl<6> vdd vss wl<3> / cell_PIM
XI17791 bl<6> cbl<3> in1<4> in2<4> sl<6> vdd vss wl<4> / cell_PIM
XI18443 bl<8> cbl<4> in1<44> in2<44> sl<8> vdd vss wl<44> / cell_PIM
XI19091 bl<20> cbl<10> in1<110> in2<110> sl<20> vdd vss wl<110> / cell_PIM
XI19090 bl<20> cbl<10> in1<109> in2<109> sl<20> vdd vss wl<109> / cell_PIM
XI19089 bl<20> cbl<10> in1<108> in2<108> sl<20> vdd vss wl<108> / cell_PIM
XI19088 bl<20> cbl<10> in1<112> in2<112> sl<20> vdd vss wl<112> / cell_PIM
XI19087 bl<20> cbl<10> in1<111> in2<111> sl<20> vdd vss wl<111> / cell_PIM
XI18437 bl<14> cbl<7> in1<49> in2<49> sl<14> vdd vss wl<49> / cell_PIM
XI18436 bl<14> cbl<7> in1<50> in2<50> sl<14> vdd vss wl<50> / cell_PIM
XI18435 bl<14> cbl<7> in1<51> in2<51> sl<14> vdd vss wl<51> / cell_PIM
XI18434 bl<14> cbl<7> in1<52> in2<52> sl<14> vdd vss wl<52> / cell_PIM
XI17786 bl<4> cbl<2> in1<4> in2<4> sl<4> vdd vss wl<4> / cell_PIM
XI17785 bl<4> cbl<2> in1<3> in2<3> sl<4> vdd vss wl<3> / cell_PIM
XI17784 bl<4> cbl<2> in1<2> in2<2> sl<4> vdd vss wl<2> / cell_PIM
XI17783 bl<4> cbl<2> in1<1> in2<1> sl<4> vdd vss wl<1> / cell_PIM
XI18433 bl<14> cbl<7> in1<48> in2<48> sl<14> vdd vss wl<48> / cell_PIM
XI19081 bl<18> cbl<9> in1<108> in2<108> sl<18> vdd vss wl<108> / cell_PIM
XI19080 bl<18> cbl<9> in1<109> in2<109> sl<18> vdd vss wl<109> / cell_PIM
XI19079 bl<18> cbl<9> in1<110> in2<110> sl<18> vdd vss wl<110> / cell_PIM
XI17777 bl<6> cbl<3> in1<6> in2<6> sl<6> vdd vss wl<6> / cell_PIM
XI17776 bl<6> cbl<3> in1<7> in2<7> sl<6> vdd vss wl<7> / cell_PIM
XI17775 bl<6> cbl<3> in1<8> in2<8> sl<6> vdd vss wl<8> / cell_PIM
XI17774 bl<6> cbl<3> in1<9> in2<9> sl<6> vdd vss wl<9> / cell_PIM
XI18427 bl<12> cbl<6> in1<52> in2<52> sl<12> vdd vss wl<52> / cell_PIM
XI18426 bl<12> cbl<6> in1<51> in2<51> sl<12> vdd vss wl<51> / cell_PIM
XI18425 bl<12> cbl<6> in1<50> in2<50> sl<12> vdd vss wl<50> / cell_PIM
XI18424 bl<12> cbl<6> in1<49> in2<49> sl<12> vdd vss wl<49> / cell_PIM
XI19078 bl<18> cbl<9> in1<112> in2<112> sl<18> vdd vss wl<112> / cell_PIM
XI19077 bl<18> cbl<9> in1<111> in2<111> sl<18> vdd vss wl<111> / cell_PIM
XI17773 bl<6> cbl<3> in1<5> in2<5> sl<6> vdd vss wl<5> / cell_PIM
XI18423 bl<12> cbl<6> in1<48> in2<48> sl<12> vdd vss wl<48> / cell_PIM
XI19071 bl<16> cbl<8> in1<110> in2<110> sl<16> vdd vss wl<110> / cell_PIM
XI19070 bl<16> cbl<8> in1<109> in2<109> sl<16> vdd vss wl<109> / cell_PIM
XI19069 bl<16> cbl<8> in1<108> in2<108> sl<16> vdd vss wl<108> / cell_PIM
XI19068 bl<16> cbl<8> in1<112> in2<112> sl<16> vdd vss wl<112> / cell_PIM
XI19067 bl<16> cbl<8> in1<111> in2<111> sl<16> vdd vss wl<111> / cell_PIM
XI18417 bl<10> cbl<5> in1<49> in2<49> sl<10> vdd vss wl<49> / cell_PIM
XI18416 bl<10> cbl<5> in1<50> in2<50> sl<10> vdd vss wl<50> / cell_PIM
XI18415 bl<10> cbl<5> in1<51> in2<51> sl<10> vdd vss wl<51> / cell_PIM
XI18414 bl<10> cbl<5> in1<52> in2<52> sl<10> vdd vss wl<52> / cell_PIM
XI17767 bl<4> cbl<2> in1<9> in2<9> sl<4> vdd vss wl<9> / cell_PIM
XI17766 bl<4> cbl<2> in1<8> in2<8> sl<4> vdd vss wl<8> / cell_PIM
XI17765 bl<4> cbl<2> in1<7> in2<7> sl<4> vdd vss wl<7> / cell_PIM
XI17764 bl<4> cbl<2> in1<6> in2<6> sl<4> vdd vss wl<6> / cell_PIM
XI17763 bl<4> cbl<2> in1<5> in2<5> sl<4> vdd vss wl<5> / cell_PIM
XI18413 bl<10> cbl<5> in1<48> in2<48> sl<10> vdd vss wl<48> / cell_PIM
XI19061 bl<30> cbl<15> in1<113> in2<113> sl<30> vdd vss wl<113> / cell_PIM
XI19060 bl<30> cbl<15> in1<114> in2<114> sl<30> vdd vss wl<114> / cell_PIM
XI19059 bl<30> cbl<15> in1<115> in2<115> sl<30> vdd vss wl<115> / cell_PIM
XI17757 bl<6> cbl<3> in1<11> in2<11> sl<6> vdd vss wl<11> / cell_PIM
XI17756 bl<6> cbl<3> in1<12> in2<12> sl<6> vdd vss wl<12> / cell_PIM
XI17755 bl<6> cbl<3> in1<13> in2<13> sl<6> vdd vss wl<13> / cell_PIM
XI17754 bl<6> cbl<3> in1<14> in2<14> sl<6> vdd vss wl<14> / cell_PIM
XI18407 bl<8> cbl<4> in1<52> in2<52> sl<8> vdd vss wl<52> / cell_PIM
XI18406 bl<8> cbl<4> in1<51> in2<51> sl<8> vdd vss wl<51> / cell_PIM
XI18405 bl<8> cbl<4> in1<50> in2<50> sl<8> vdd vss wl<50> / cell_PIM
XI18404 bl<8> cbl<4> in1<49> in2<49> sl<8> vdd vss wl<49> / cell_PIM
XI19058 bl<30> cbl<15> in1<117> in2<117> sl<30> vdd vss wl<117> / cell_PIM
XI19057 bl<30> cbl<15> in1<116> in2<116> sl<30> vdd vss wl<116> / cell_PIM
XI17753 bl<6> cbl<3> in1<10> in2<10> sl<6> vdd vss wl<10> / cell_PIM
XI18403 bl<8> cbl<4> in1<48> in2<48> sl<8> vdd vss wl<48> / cell_PIM
XI19051 bl<28> cbl<14> in1<115> in2<115> sl<28> vdd vss wl<115> / cell_PIM
XI19050 bl<28> cbl<14> in1<114> in2<114> sl<28> vdd vss wl<114> / cell_PIM
XI19049 bl<28> cbl<14> in1<113> in2<113> sl<28> vdd vss wl<113> / cell_PIM
XI19048 bl<28> cbl<14> in1<117> in2<117> sl<28> vdd vss wl<117> / cell_PIM
XI19047 bl<28> cbl<14> in1<116> in2<116> sl<28> vdd vss wl<116> / cell_PIM
XI18397 bl<14> cbl<7> in1<54> in2<54> sl<14> vdd vss wl<54> / cell_PIM
XI18396 bl<14> cbl<7> in1<55> in2<55> sl<14> vdd vss wl<55> / cell_PIM
XI18395 bl<14> cbl<7> in1<56> in2<56> sl<14> vdd vss wl<56> / cell_PIM
XI18394 bl<14> cbl<7> in1<57> in2<57> sl<14> vdd vss wl<57> / cell_PIM
XI17747 bl<4> cbl<2> in1<14> in2<14> sl<4> vdd vss wl<14> / cell_PIM
XI17746 bl<4> cbl<2> in1<13> in2<13> sl<4> vdd vss wl<13> / cell_PIM
XI17745 bl<4> cbl<2> in1<12> in2<12> sl<4> vdd vss wl<12> / cell_PIM
XI17744 bl<4> cbl<2> in1<11> in2<11> sl<4> vdd vss wl<11> / cell_PIM
XI17743 bl<4> cbl<2> in1<10> in2<10> sl<4> vdd vss wl<10> / cell_PIM
XI18393 bl<14> cbl<7> in1<53> in2<53> sl<14> vdd vss wl<53> / cell_PIM
XI19041 bl<26> cbl<13> in1<113> in2<113> sl<26> vdd vss wl<113> / cell_PIM
XI19040 bl<26> cbl<13> in1<114> in2<114> sl<26> vdd vss wl<114> / cell_PIM
XI19039 bl<26> cbl<13> in1<115> in2<115> sl<26> vdd vss wl<115> / cell_PIM
XI17737 bl<6> cbl<3> in1<16> in2<16> sl<6> vdd vss wl<16> / cell_PIM
XI17736 bl<6> cbl<3> in1<17> in2<17> sl<6> vdd vss wl<17> / cell_PIM
XI17735 bl<6> cbl<3> in1<18> in2<18> sl<6> vdd vss wl<18> / cell_PIM
XI17734 bl<6> cbl<3> in1<19> in2<19> sl<6> vdd vss wl<19> / cell_PIM
XI18387 bl<12> cbl<6> in1<57> in2<57> sl<12> vdd vss wl<57> / cell_PIM
XI18386 bl<12> cbl<6> in1<56> in2<56> sl<12> vdd vss wl<56> / cell_PIM
XI18385 bl<12> cbl<6> in1<55> in2<55> sl<12> vdd vss wl<55> / cell_PIM
XI18384 bl<12> cbl<6> in1<54> in2<54> sl<12> vdd vss wl<54> / cell_PIM
XI19038 bl<26> cbl<13> in1<117> in2<117> sl<26> vdd vss wl<117> / cell_PIM
XI19037 bl<26> cbl<13> in1<116> in2<116> sl<26> vdd vss wl<116> / cell_PIM
XI17733 bl<6> cbl<3> in1<15> in2<15> sl<6> vdd vss wl<15> / cell_PIM
XI18383 bl<12> cbl<6> in1<53> in2<53> sl<12> vdd vss wl<53> / cell_PIM
XI19031 bl<24> cbl<12> in1<113> in2<113> sl<24> vdd vss wl<113> / cell_PIM
XI19030 bl<24> cbl<12> in1<114> in2<114> sl<24> vdd vss wl<114> / cell_PIM
XI19029 bl<24> cbl<12> in1<115> in2<115> sl<24> vdd vss wl<115> / cell_PIM
XI19028 bl<24> cbl<12> in1<117> in2<117> sl<24> vdd vss wl<117> / cell_PIM
XI19027 bl<24> cbl<12> in1<116> in2<116> sl<24> vdd vss wl<116> / cell_PIM
XI18377 bl<10> cbl<5> in1<54> in2<54> sl<10> vdd vss wl<54> / cell_PIM
XI18376 bl<10> cbl<5> in1<55> in2<55> sl<10> vdd vss wl<55> / cell_PIM
XI18375 bl<10> cbl<5> in1<56> in2<56> sl<10> vdd vss wl<56> / cell_PIM
XI18374 bl<10> cbl<5> in1<57> in2<57> sl<10> vdd vss wl<57> / cell_PIM
XI17727 bl<4> cbl<2> in1<19> in2<19> sl<4> vdd vss wl<19> / cell_PIM
XI17726 bl<4> cbl<2> in1<18> in2<18> sl<4> vdd vss wl<18> / cell_PIM
XI17725 bl<4> cbl<2> in1<17> in2<17> sl<4> vdd vss wl<17> / cell_PIM
XI17724 bl<4> cbl<2> in1<16> in2<16> sl<4> vdd vss wl<16> / cell_PIM
XI17723 bl<4> cbl<2> in1<15> in2<15> sl<4> vdd vss wl<15> / cell_PIM
XI18373 bl<10> cbl<5> in1<53> in2<53> sl<10> vdd vss wl<53> / cell_PIM
XI19021 bl<22> cbl<11> in1<113> in2<113> sl<22> vdd vss wl<113> / cell_PIM
XI19020 bl<22> cbl<11> in1<114> in2<114> sl<22> vdd vss wl<114> / cell_PIM
XI19019 bl<22> cbl<11> in1<115> in2<115> sl<22> vdd vss wl<115> / cell_PIM
XI17717 bl<6> cbl<3> in1<21> in2<21> sl<6> vdd vss wl<21> / cell_PIM
XI17716 bl<6> cbl<3> in1<22> in2<22> sl<6> vdd vss wl<22> / cell_PIM
XI17715 bl<6> cbl<3> in1<23> in2<23> sl<6> vdd vss wl<23> / cell_PIM
XI17714 bl<6> cbl<3> in1<24> in2<24> sl<6> vdd vss wl<24> / cell_PIM
XI18367 bl<8> cbl<4> in1<57> in2<57> sl<8> vdd vss wl<57> / cell_PIM
XI18366 bl<8> cbl<4> in1<56> in2<56> sl<8> vdd vss wl<56> / cell_PIM
XI18365 bl<8> cbl<4> in1<55> in2<55> sl<8> vdd vss wl<55> / cell_PIM
XI18364 bl<8> cbl<4> in1<54> in2<54> sl<8> vdd vss wl<54> / cell_PIM
XI19018 bl<22> cbl<11> in1<117> in2<117> sl<22> vdd vss wl<117> / cell_PIM
XI19017 bl<22> cbl<11> in1<116> in2<116> sl<22> vdd vss wl<116> / cell_PIM
XI17713 bl<6> cbl<3> in1<20> in2<20> sl<6> vdd vss wl<20> / cell_PIM
XI18363 bl<8> cbl<4> in1<53> in2<53> sl<8> vdd vss wl<53> / cell_PIM
XI19011 bl<20> cbl<10> in1<115> in2<115> sl<20> vdd vss wl<115> / cell_PIM
XI19010 bl<20> cbl<10> in1<114> in2<114> sl<20> vdd vss wl<114> / cell_PIM
XI19009 bl<20> cbl<10> in1<113> in2<113> sl<20> vdd vss wl<113> / cell_PIM
XI19008 bl<20> cbl<10> in1<117> in2<117> sl<20> vdd vss wl<117> / cell_PIM
XI19007 bl<20> cbl<10> in1<116> in2<116> sl<20> vdd vss wl<116> / cell_PIM
XI18357 bl<14> cbl<7> in1<59> in2<59> sl<14> vdd vss wl<59> / cell_PIM
XI18356 bl<14> cbl<7> in1<60> in2<60> sl<14> vdd vss wl<60> / cell_PIM
XI18355 bl<14> cbl<7> in1<61> in2<61> sl<14> vdd vss wl<61> / cell_PIM
XI18354 bl<14> cbl<7> in1<62> in2<62> sl<14> vdd vss wl<62> / cell_PIM
XI17707 bl<4> cbl<2> in1<24> in2<24> sl<4> vdd vss wl<24> / cell_PIM
XI17706 bl<4> cbl<2> in1<23> in2<23> sl<4> vdd vss wl<23> / cell_PIM
XI17705 bl<4> cbl<2> in1<22> in2<22> sl<4> vdd vss wl<22> / cell_PIM
XI17704 bl<4> cbl<2> in1<21> in2<21> sl<4> vdd vss wl<21> / cell_PIM
XI17703 bl<4> cbl<2> in1<20> in2<20> sl<4> vdd vss wl<20> / cell_PIM
XI18353 bl<14> cbl<7> in1<58> in2<58> sl<14> vdd vss wl<58> / cell_PIM
XI19001 bl<18> cbl<9> in1<113> in2<113> sl<18> vdd vss wl<113> / cell_PIM
XI19000 bl<18> cbl<9> in1<114> in2<114> sl<18> vdd vss wl<114> / cell_PIM
XI18999 bl<18> cbl<9> in1<115> in2<115> sl<18> vdd vss wl<115> / cell_PIM
XI17698 bl<6> cbl<3> in1<26> in2<26> sl<6> vdd vss wl<26> / cell_PIM
XI17697 bl<6> cbl<3> in1<27> in2<27> sl<6> vdd vss wl<27> / cell_PIM
XI17696 bl<6> cbl<3> in1<28> in2<28> sl<6> vdd vss wl<28> / cell_PIM
XI17695 bl<6> cbl<3> in1<25> in2<25> sl<6> vdd vss wl<25> / cell_PIM
XI18347 bl<12> cbl<6> in1<62> in2<62> sl<12> vdd vss wl<62> / cell_PIM
XI18346 bl<12> cbl<6> in1<61> in2<61> sl<12> vdd vss wl<61> / cell_PIM
XI18345 bl<12> cbl<6> in1<60> in2<60> sl<12> vdd vss wl<60> / cell_PIM
XI18344 bl<12> cbl<6> in1<59> in2<59> sl<12> vdd vss wl<59> / cell_PIM
XI18998 bl<18> cbl<9> in1<117> in2<117> sl<18> vdd vss wl<117> / cell_PIM
XI18997 bl<18> cbl<9> in1<116> in2<116> sl<18> vdd vss wl<116> / cell_PIM
XI17690 bl<4> cbl<2> in1<28> in2<28> sl<4> vdd vss wl<28> / cell_PIM
XI17689 bl<4> cbl<2> in1<27> in2<27> sl<4> vdd vss wl<27> / cell_PIM
XI18343 bl<12> cbl<6> in1<58> in2<58> sl<12> vdd vss wl<58> / cell_PIM
XI18991 bl<16> cbl<8> in1<115> in2<115> sl<16> vdd vss wl<115> / cell_PIM
XI18990 bl<16> cbl<8> in1<114> in2<114> sl<16> vdd vss wl<114> / cell_PIM
XI18989 bl<16> cbl<8> in1<113> in2<113> sl<16> vdd vss wl<113> / cell_PIM
XI18988 bl<16> cbl<8> in1<117> in2<117> sl<16> vdd vss wl<117> / cell_PIM
XI18987 bl<16> cbl<8> in1<116> in2<116> sl<16> vdd vss wl<116> / cell_PIM
XI18337 bl<10> cbl<5> in1<59> in2<59> sl<10> vdd vss wl<59> / cell_PIM
XI18336 bl<10> cbl<5> in1<60> in2<60> sl<10> vdd vss wl<60> / cell_PIM
XI18335 bl<10> cbl<5> in1<61> in2<61> sl<10> vdd vss wl<61> / cell_PIM
XI18334 bl<10> cbl<5> in1<62> in2<62> sl<10> vdd vss wl<62> / cell_PIM
XI17688 bl<4> cbl<2> in1<26> in2<26> sl<4> vdd vss wl<26> / cell_PIM
XI17687 bl<4> cbl<2> in1<25> in2<25> sl<4> vdd vss wl<25> / cell_PIM
XI17681 bl<6> cbl<3> in1<30> in2<30> sl<6> vdd vss wl<30> / cell_PIM
XI17680 bl<6> cbl<3> in1<31> in2<31> sl<6> vdd vss wl<31> / cell_PIM
XI17679 bl<6> cbl<3> in1<32> in2<32> sl<6> vdd vss wl<32> / cell_PIM
XI18333 bl<10> cbl<5> in1<58> in2<58> sl<10> vdd vss wl<58> / cell_PIM
XI18981 bl<30> cbl<15> in1<118> in2<118> sl<30> vdd vss wl<118> / cell_PIM
XI18980 bl<30> cbl<15> in1<119> in2<119> sl<30> vdd vss wl<119> / cell_PIM
XI18979 bl<30> cbl<15> in1<121> in2<121> sl<30> vdd vss wl<121> / cell_PIM
XI17678 bl<6> cbl<3> in1<33> in2<33> sl<6> vdd vss wl<33> / cell_PIM
XI17677 bl<6> cbl<3> in1<29> in2<29> sl<6> vdd vss wl<29> / cell_PIM
XI18327 bl<8> cbl<4> in1<62> in2<62> sl<8> vdd vss wl<62> / cell_PIM
XI18326 bl<8> cbl<4> in1<61> in2<61> sl<8> vdd vss wl<61> / cell_PIM
XI18325 bl<8> cbl<4> in1<60> in2<60> sl<8> vdd vss wl<60> / cell_PIM
XI18324 bl<8> cbl<4> in1<59> in2<59> sl<8> vdd vss wl<59> / cell_PIM
XI18978 bl<30> cbl<15> in1<122> in2<122> sl<30> vdd vss wl<122> / cell_PIM
XI18977 bl<30> cbl<15> in1<120> in2<120> sl<30> vdd vss wl<120> / cell_PIM
XI17671 bl<4> cbl<2> in1<33> in2<33> sl<4> vdd vss wl<33> / cell_PIM
XI17670 bl<4> cbl<2> in1<32> in2<32> sl<4> vdd vss wl<32> / cell_PIM
XI17669 bl<4> cbl<2> in1<31> in2<31> sl<4> vdd vss wl<31> / cell_PIM
XI18323 bl<8> cbl<4> in1<58> in2<58> sl<8> vdd vss wl<58> / cell_PIM
XI18971 bl<28> cbl<14> in1<119> in2<119> sl<28> vdd vss wl<119> / cell_PIM
XI18970 bl<28> cbl<14> in1<118> in2<118> sl<28> vdd vss wl<118> / cell_PIM
XI18969 bl<28> cbl<14> in1<122> in2<122> sl<28> vdd vss wl<122> / cell_PIM
XI18968 bl<28> cbl<14> in1<121> in2<121> sl<28> vdd vss wl<121> / cell_PIM
XI18967 bl<28> cbl<14> in1<120> in2<120> sl<28> vdd vss wl<120> / cell_PIM
XI18317 bl<14> cbl<7> in1<64> in2<64> sl<14> vdd vss wl<64> / cell_PIM
XI18316 bl<14> cbl<7> in1<65> in2<65> sl<14> vdd vss wl<65> / cell_PIM
XI18315 bl<14> cbl<7> in1<66> in2<66> sl<14> vdd vss wl<66> / cell_PIM
XI18314 bl<14> cbl<7> in1<67> in2<67> sl<14> vdd vss wl<67> / cell_PIM
XI17668 bl<4> cbl<2> in1<30> in2<30> sl<4> vdd vss wl<30> / cell_PIM
XI17667 bl<4> cbl<2> in1<29> in2<29> sl<4> vdd vss wl<29> / cell_PIM
XI17661 bl<6> cbl<3> in1<35> in2<35> sl<6> vdd vss wl<35> / cell_PIM
XI17660 bl<6> cbl<3> in1<36> in2<36> sl<6> vdd vss wl<36> / cell_PIM
XI17659 bl<6> cbl<3> in1<37> in2<37> sl<6> vdd vss wl<37> / cell_PIM
XI18313 bl<14> cbl<7> in1<63> in2<63> sl<14> vdd vss wl<63> / cell_PIM
XI18961 bl<26> cbl<13> in1<118> in2<118> sl<26> vdd vss wl<118> / cell_PIM
XI18960 bl<26> cbl<13> in1<119> in2<119> sl<26> vdd vss wl<119> / cell_PIM
XI18959 bl<26> cbl<13> in1<121> in2<121> sl<26> vdd vss wl<121> / cell_PIM
XI17658 bl<6> cbl<3> in1<38> in2<38> sl<6> vdd vss wl<38> / cell_PIM
XI17657 bl<6> cbl<3> in1<34> in2<34> sl<6> vdd vss wl<34> / cell_PIM
XI18307 bl<12> cbl<6> in1<67> in2<67> sl<12> vdd vss wl<67> / cell_PIM
XI18306 bl<12> cbl<6> in1<66> in2<66> sl<12> vdd vss wl<66> / cell_PIM
XI18305 bl<12> cbl<6> in1<65> in2<65> sl<12> vdd vss wl<65> / cell_PIM
XI18304 bl<12> cbl<6> in1<64> in2<64> sl<12> vdd vss wl<64> / cell_PIM
XI18958 bl<26> cbl<13> in1<122> in2<122> sl<26> vdd vss wl<122> / cell_PIM
XI18957 bl<26> cbl<13> in1<120> in2<120> sl<26> vdd vss wl<120> / cell_PIM
XI17651 bl<4> cbl<2> in1<38> in2<38> sl<4> vdd vss wl<38> / cell_PIM
XI17650 bl<4> cbl<2> in1<37> in2<37> sl<4> vdd vss wl<37> / cell_PIM
XI17649 bl<4> cbl<2> in1<36> in2<36> sl<4> vdd vss wl<36> / cell_PIM
XI18303 bl<12> cbl<6> in1<63> in2<63> sl<12> vdd vss wl<63> / cell_PIM
XI18951 bl<24> cbl<12> in1<118> in2<118> sl<24> vdd vss wl<118> / cell_PIM
XI18950 bl<24> cbl<12> in1<119> in2<119> sl<24> vdd vss wl<119> / cell_PIM
XI18949 bl<24> cbl<12> in1<121> in2<121> sl<24> vdd vss wl<121> / cell_PIM
XI18948 bl<24> cbl<12> in1<122> in2<122> sl<24> vdd vss wl<122> / cell_PIM
XI18947 bl<24> cbl<12> in1<120> in2<120> sl<24> vdd vss wl<120> / cell_PIM
XI18297 bl<10> cbl<5> in1<64> in2<64> sl<10> vdd vss wl<64> / cell_PIM
XI18296 bl<10> cbl<5> in1<65> in2<65> sl<10> vdd vss wl<65> / cell_PIM
XI18295 bl<10> cbl<5> in1<66> in2<66> sl<10> vdd vss wl<66> / cell_PIM
XI18294 bl<10> cbl<5> in1<67> in2<67> sl<10> vdd vss wl<67> / cell_PIM
XI17648 bl<4> cbl<2> in1<35> in2<35> sl<4> vdd vss wl<35> / cell_PIM
XI17647 bl<4> cbl<2> in1<34> in2<34> sl<4> vdd vss wl<34> / cell_PIM
XI17641 bl<6> cbl<3> in1<40> in2<40> sl<6> vdd vss wl<40> / cell_PIM
XI17640 bl<6> cbl<3> in1<41> in2<41> sl<6> vdd vss wl<41> / cell_PIM
XI17639 bl<6> cbl<3> in1<42> in2<42> sl<6> vdd vss wl<42> / cell_PIM
XI18293 bl<10> cbl<5> in1<63> in2<63> sl<10> vdd vss wl<63> / cell_PIM
XI18941 bl<22> cbl<11> in1<118> in2<118> sl<22> vdd vss wl<118> / cell_PIM
XI18940 bl<22> cbl<11> in1<119> in2<119> sl<22> vdd vss wl<119> / cell_PIM
XI18939 bl<22> cbl<11> in1<121> in2<121> sl<22> vdd vss wl<121> / cell_PIM
XI17638 bl<6> cbl<3> in1<43> in2<43> sl<6> vdd vss wl<43> / cell_PIM
XI17637 bl<6> cbl<3> in1<39> in2<39> sl<6> vdd vss wl<39> / cell_PIM
XI18287 bl<8> cbl<4> in1<67> in2<67> sl<8> vdd vss wl<67> / cell_PIM
XI18286 bl<8> cbl<4> in1<66> in2<66> sl<8> vdd vss wl<66> / cell_PIM
XI18285 bl<8> cbl<4> in1<65> in2<65> sl<8> vdd vss wl<65> / cell_PIM
XI18284 bl<8> cbl<4> in1<64> in2<64> sl<8> vdd vss wl<64> / cell_PIM
XI18938 bl<22> cbl<11> in1<122> in2<122> sl<22> vdd vss wl<122> / cell_PIM
XI18937 bl<22> cbl<11> in1<120> in2<120> sl<22> vdd vss wl<120> / cell_PIM
XI17631 bl<4> cbl<2> in1<43> in2<43> sl<4> vdd vss wl<43> / cell_PIM
XI17630 bl<4> cbl<2> in1<42> in2<42> sl<4> vdd vss wl<42> / cell_PIM
XI17629 bl<4> cbl<2> in1<41> in2<41> sl<4> vdd vss wl<41> / cell_PIM
XI18283 bl<8> cbl<4> in1<63> in2<63> sl<8> vdd vss wl<63> / cell_PIM
XI18931 bl<20> cbl<10> in1<119> in2<119> sl<20> vdd vss wl<119> / cell_PIM
XI18930 bl<20> cbl<10> in1<118> in2<118> sl<20> vdd vss wl<118> / cell_PIM
XI18929 bl<20> cbl<10> in1<122> in2<122> sl<20> vdd vss wl<122> / cell_PIM
XI18928 bl<20> cbl<10> in1<121> in2<121> sl<20> vdd vss wl<121> / cell_PIM
XI18927 bl<20> cbl<10> in1<120> in2<120> sl<20> vdd vss wl<120> / cell_PIM
XI18278 bl<14> cbl<7> in1<69> in2<69> sl<14> vdd vss wl<69> / cell_PIM
XI18277 bl<14> cbl<7> in1<70> in2<70> sl<14> vdd vss wl<70> / cell_PIM
XI18276 bl<14> cbl<7> in1<71> in2<71> sl<14> vdd vss wl<71> / cell_PIM
XI18275 bl<14> cbl<7> in1<68> in2<68> sl<14> vdd vss wl<68> / cell_PIM
XI17628 bl<4> cbl<2> in1<40> in2<40> sl<4> vdd vss wl<40> / cell_PIM
XI17627 bl<4> cbl<2> in1<39> in2<39> sl<4> vdd vss wl<39> / cell_PIM
XI17622 bl<6> cbl<3> in1<45> in2<45> sl<6> vdd vss wl<45> / cell_PIM
XI17621 bl<6> cbl<3> in1<46> in2<46> sl<6> vdd vss wl<46> / cell_PIM
XI17620 bl<6> cbl<3> in1<47> in2<47> sl<6> vdd vss wl<47> / cell_PIM
XI17619 bl<6> cbl<3> in1<44> in2<44> sl<6> vdd vss wl<44> / cell_PIM
XI18270 bl<12> cbl<6> in1<71> in2<71> sl<12> vdd vss wl<71> / cell_PIM
XI18269 bl<12> cbl<6> in1<70> in2<70> sl<12> vdd vss wl<70> / cell_PIM
XI18921 bl<18> cbl<9> in1<118> in2<118> sl<18> vdd vss wl<118> / cell_PIM
XI18920 bl<18> cbl<9> in1<119> in2<119> sl<18> vdd vss wl<119> / cell_PIM
XI18919 bl<18> cbl<9> in1<121> in2<121> sl<18> vdd vss wl<121> / cell_PIM
XI17614 bl<4> cbl<2> in1<47> in2<47> sl<4> vdd vss wl<47> / cell_PIM
XI18268 bl<12> cbl<6> in1<69> in2<69> sl<12> vdd vss wl<69> / cell_PIM
XI18267 bl<12> cbl<6> in1<68> in2<68> sl<12> vdd vss wl<68> / cell_PIM
XI18918 bl<18> cbl<9> in1<122> in2<122> sl<18> vdd vss wl<122> / cell_PIM
XI18917 bl<18> cbl<9> in1<120> in2<120> sl<18> vdd vss wl<120> / cell_PIM
XI17613 bl<4> cbl<2> in1<46> in2<46> sl<4> vdd vss wl<46> / cell_PIM
XI17612 bl<4> cbl<2> in1<45> in2<45> sl<4> vdd vss wl<45> / cell_PIM
XI17611 bl<4> cbl<2> in1<44> in2<44> sl<4> vdd vss wl<44> / cell_PIM
XI18262 bl<10> cbl<5> in1<69> in2<69> sl<10> vdd vss wl<69> / cell_PIM
XI18261 bl<10> cbl<5> in1<70> in2<70> sl<10> vdd vss wl<70> / cell_PIM
XI18260 bl<10> cbl<5> in1<71> in2<71> sl<10> vdd vss wl<71> / cell_PIM
XI18259 bl<10> cbl<5> in1<68> in2<68> sl<10> vdd vss wl<68> / cell_PIM
XI18911 bl<16> cbl<8> in1<119> in2<119> sl<16> vdd vss wl<119> / cell_PIM
XI18910 bl<16> cbl<8> in1<118> in2<118> sl<16> vdd vss wl<118> / cell_PIM
XI18909 bl<16> cbl<8> in1<122> in2<122> sl<16> vdd vss wl<122> / cell_PIM
XI18908 bl<16> cbl<8> in1<121> in2<121> sl<16> vdd vss wl<121> / cell_PIM
XI18907 bl<16> cbl<8> in1<120> in2<120> sl<16> vdd vss wl<120> / cell_PIM
XI18254 bl<8> cbl<4> in1<71> in2<71> sl<8> vdd vss wl<71> / cell_PIM
XI17605 bl<6> cbl<3> in1<49> in2<49> sl<6> vdd vss wl<49> / cell_PIM
XI17604 bl<6> cbl<3> in1<50> in2<50> sl<6> vdd vss wl<50> / cell_PIM
XI17603 bl<6> cbl<3> in1<51> in2<51> sl<6> vdd vss wl<51> / cell_PIM
XI17602 bl<6> cbl<3> in1<52> in2<52> sl<6> vdd vss wl<52> / cell_PIM
XI17601 bl<6> cbl<3> in1<48> in2<48> sl<6> vdd vss wl<48> / cell_PIM
XI18253 bl<8> cbl<4> in1<70> in2<70> sl<8> vdd vss wl<70> / cell_PIM
XI18252 bl<8> cbl<4> in1<69> in2<69> sl<8> vdd vss wl<69> / cell_PIM
XI18251 bl<8> cbl<4> in1<68> in2<68> sl<8> vdd vss wl<68> / cell_PIM
XI18901 bl<30> cbl<15> in1<127> in2<127> sl<30> vdd vss wl<127> / cell_PIM
XI18900 bl<30> cbl<15> in1<126> in2<126> sl<30> vdd vss wl<126> / cell_PIM
XI18899 bl<30> cbl<15> in1<125> in2<125> sl<30> vdd vss wl<125> / cell_PIM
XI17595 bl<4> cbl<2> in1<52> in2<52> sl<4> vdd vss wl<52> / cell_PIM
XI17594 bl<4> cbl<2> in1<51> in2<51> sl<4> vdd vss wl<51> / cell_PIM
XI18245 bl<14> cbl<7> in1<73> in2<73> sl<14> vdd vss wl<73> / cell_PIM
XI18244 bl<14> cbl<7> in1<74> in2<74> sl<14> vdd vss wl<74> / cell_PIM
XI18898 bl<30> cbl<15> in1<123> in2<123> sl<30> vdd vss wl<123> / cell_PIM
XI18897 bl<30> cbl<15> in1<124> in2<124> sl<30> vdd vss wl<124> / cell_PIM
XI17593 bl<4> cbl<2> in1<50> in2<50> sl<4> vdd vss wl<50> / cell_PIM
XI17592 bl<4> cbl<2> in1<49> in2<49> sl<4> vdd vss wl<49> / cell_PIM
XI17591 bl<4> cbl<2> in1<48> in2<48> sl<4> vdd vss wl<48> / cell_PIM
XI18243 bl<14> cbl<7> in1<75> in2<75> sl<14> vdd vss wl<75> / cell_PIM
XI18242 bl<14> cbl<7> in1<76> in2<76> sl<14> vdd vss wl<76> / cell_PIM
XI18241 bl<14> cbl<7> in1<72> in2<72> sl<14> vdd vss wl<72> / cell_PIM
XI18891 bl<28> cbl<14> in1<127> in2<127> sl<28> vdd vss wl<127> / cell_PIM
XI18890 bl<28> cbl<14> in1<126> in2<126> sl<28> vdd vss wl<126> / cell_PIM
XI18889 bl<28> cbl<14> in1<125> in2<125> sl<28> vdd vss wl<125> / cell_PIM
XI18888 bl<28> cbl<14> in1<124> in2<124> sl<28> vdd vss wl<124> / cell_PIM
XI18887 bl<28> cbl<14> in1<123> in2<123> sl<28> vdd vss wl<123> / cell_PIM
XI18235 bl<12> cbl<6> in1<76> in2<76> sl<12> vdd vss wl<76> / cell_PIM
XI18234 bl<12> cbl<6> in1<75> in2<75> sl<12> vdd vss wl<75> / cell_PIM
XI17585 bl<6> cbl<3> in1<54> in2<54> sl<6> vdd vss wl<54> / cell_PIM
XI17584 bl<6> cbl<3> in1<55> in2<55> sl<6> vdd vss wl<55> / cell_PIM
XI17583 bl<6> cbl<3> in1<56> in2<56> sl<6> vdd vss wl<56> / cell_PIM
XI17582 bl<6> cbl<3> in1<57> in2<57> sl<6> vdd vss wl<57> / cell_PIM
XI17581 bl<6> cbl<3> in1<53> in2<53> sl<6> vdd vss wl<53> / cell_PIM
XI18233 bl<12> cbl<6> in1<74> in2<74> sl<12> vdd vss wl<74> / cell_PIM
XI18232 bl<12> cbl<6> in1<73> in2<73> sl<12> vdd vss wl<73> / cell_PIM
XI18231 bl<12> cbl<6> in1<72> in2<72> sl<12> vdd vss wl<72> / cell_PIM
XI18881 bl<26> cbl<13> in1<127> in2<127> sl<26> vdd vss wl<127> / cell_PIM
XI18880 bl<26> cbl<13> in1<126> in2<126> sl<26> vdd vss wl<126> / cell_PIM
XI18879 bl<26> cbl<13> in1<125> in2<125> sl<26> vdd vss wl<125> / cell_PIM
XI17575 bl<4> cbl<2> in1<57> in2<57> sl<4> vdd vss wl<57> / cell_PIM
XI17574 bl<4> cbl<2> in1<56> in2<56> sl<4> vdd vss wl<56> / cell_PIM
XI18225 bl<10> cbl<5> in1<73> in2<73> sl<10> vdd vss wl<73> / cell_PIM
XI18224 bl<10> cbl<5> in1<74> in2<74> sl<10> vdd vss wl<74> / cell_PIM
XI18878 bl<26> cbl<13> in1<123> in2<123> sl<26> vdd vss wl<123> / cell_PIM
XI18877 bl<26> cbl<13> in1<124> in2<124> sl<26> vdd vss wl<124> / cell_PIM
XI17573 bl<4> cbl<2> in1<55> in2<55> sl<4> vdd vss wl<55> / cell_PIM
XI17572 bl<4> cbl<2> in1<54> in2<54> sl<4> vdd vss wl<54> / cell_PIM
XI17571 bl<4> cbl<2> in1<53> in2<53> sl<4> vdd vss wl<53> / cell_PIM
XI18223 bl<10> cbl<5> in1<75> in2<75> sl<10> vdd vss wl<75> / cell_PIM
XI18222 bl<10> cbl<5> in1<76> in2<76> sl<10> vdd vss wl<76> / cell_PIM
XI18221 bl<10> cbl<5> in1<72> in2<72> sl<10> vdd vss wl<72> / cell_PIM
XI18871 bl<24> cbl<12> in1<127> in2<127> sl<24> vdd vss wl<127> / cell_PIM
XI18870 bl<24> cbl<12> in1<126> in2<126> sl<24> vdd vss wl<126> / cell_PIM
XI18869 bl<24> cbl<12> in1<125> in2<125> sl<24> vdd vss wl<125> / cell_PIM
XI18868 bl<24> cbl<12> in1<123> in2<123> sl<24> vdd vss wl<123> / cell_PIM
XI18867 bl<24> cbl<12> in1<124> in2<124> sl<24> vdd vss wl<124> / cell_PIM
XI18215 bl<8> cbl<4> in1<76> in2<76> sl<8> vdd vss wl<76> / cell_PIM
XI18214 bl<8> cbl<4> in1<75> in2<75> sl<8> vdd vss wl<75> / cell_PIM
XI17565 bl<6> cbl<3> in1<59> in2<59> sl<6> vdd vss wl<59> / cell_PIM
XI17564 bl<6> cbl<3> in1<60> in2<60> sl<6> vdd vss wl<60> / cell_PIM
XI17563 bl<6> cbl<3> in1<61> in2<61> sl<6> vdd vss wl<61> / cell_PIM
XI17562 bl<6> cbl<3> in1<62> in2<62> sl<6> vdd vss wl<62> / cell_PIM
XI17561 bl<6> cbl<3> in1<58> in2<58> sl<6> vdd vss wl<58> / cell_PIM
XI18213 bl<8> cbl<4> in1<74> in2<74> sl<8> vdd vss wl<74> / cell_PIM
XI18212 bl<8> cbl<4> in1<73> in2<73> sl<8> vdd vss wl<73> / cell_PIM
XI18211 bl<8> cbl<4> in1<72> in2<72> sl<8> vdd vss wl<72> / cell_PIM
XI18861 bl<22> cbl<11> in1<127> in2<127> sl<22> vdd vss wl<127> / cell_PIM
XI18860 bl<22> cbl<11> in1<126> in2<126> sl<22> vdd vss wl<126> / cell_PIM
XI18859 bl<22> cbl<11> in1<125> in2<125> sl<22> vdd vss wl<125> / cell_PIM
XI17555 bl<4> cbl<2> in1<62> in2<62> sl<4> vdd vss wl<62> / cell_PIM
XI17554 bl<4> cbl<2> in1<61> in2<61> sl<4> vdd vss wl<61> / cell_PIM
XI18205 bl<14> cbl<7> in1<78> in2<78> sl<14> vdd vss wl<78> / cell_PIM
XI18204 bl<14> cbl<7> in1<79> in2<79> sl<14> vdd vss wl<79> / cell_PIM
XI18858 bl<22> cbl<11> in1<123> in2<123> sl<22> vdd vss wl<123> / cell_PIM
XI18857 bl<22> cbl<11> in1<124> in2<124> sl<22> vdd vss wl<124> / cell_PIM
XI17553 bl<4> cbl<2> in1<60> in2<60> sl<4> vdd vss wl<60> / cell_PIM
XI17552 bl<4> cbl<2> in1<59> in2<59> sl<4> vdd vss wl<59> / cell_PIM
XI17551 bl<4> cbl<2> in1<58> in2<58> sl<4> vdd vss wl<58> / cell_PIM
XI18203 bl<14> cbl<7> in1<80> in2<80> sl<14> vdd vss wl<80> / cell_PIM
XI18202 bl<14> cbl<7> in1<81> in2<81> sl<14> vdd vss wl<81> / cell_PIM
XI18201 bl<14> cbl<7> in1<77> in2<77> sl<14> vdd vss wl<77> / cell_PIM
XI18851 bl<20> cbl<10> in1<127> in2<127> sl<20> vdd vss wl<127> / cell_PIM
XI18850 bl<20> cbl<10> in1<126> in2<126> sl<20> vdd vss wl<126> / cell_PIM
XI18849 bl<20> cbl<10> in1<125> in2<125> sl<20> vdd vss wl<125> / cell_PIM
XI18848 bl<20> cbl<10> in1<124> in2<124> sl<20> vdd vss wl<124> / cell_PIM
XI18847 bl<20> cbl<10> in1<123> in2<123> sl<20> vdd vss wl<123> / cell_PIM
XI18195 bl<12> cbl<6> in1<81> in2<81> sl<12> vdd vss wl<81> / cell_PIM
XI18194 bl<12> cbl<6> in1<80> in2<80> sl<12> vdd vss wl<80> / cell_PIM
XI17545 bl<6> cbl<3> in1<64> in2<64> sl<6> vdd vss wl<64> / cell_PIM
XI17544 bl<6> cbl<3> in1<65> in2<65> sl<6> vdd vss wl<65> / cell_PIM
XI17543 bl<6> cbl<3> in1<66> in2<66> sl<6> vdd vss wl<66> / cell_PIM
XI17542 bl<6> cbl<3> in1<67> in2<67> sl<6> vdd vss wl<67> / cell_PIM
XI17541 bl<6> cbl<3> in1<63> in2<63> sl<6> vdd vss wl<63> / cell_PIM
XI18193 bl<12> cbl<6> in1<79> in2<79> sl<12> vdd vss wl<79> / cell_PIM
XI18192 bl<12> cbl<6> in1<78> in2<78> sl<12> vdd vss wl<78> / cell_PIM
XI18191 bl<12> cbl<6> in1<77> in2<77> sl<12> vdd vss wl<77> / cell_PIM
XI18841 bl<18> cbl<9> in1<127> in2<127> sl<18> vdd vss wl<127> / cell_PIM
XI18840 bl<18> cbl<9> in1<126> in2<126> sl<18> vdd vss wl<126> / cell_PIM
XI18839 bl<18> cbl<9> in1<125> in2<125> sl<18> vdd vss wl<125> / cell_PIM
XI17535 bl<4> cbl<2> in1<67> in2<67> sl<4> vdd vss wl<67> / cell_PIM
XI17534 bl<4> cbl<2> in1<66> in2<66> sl<4> vdd vss wl<66> / cell_PIM
XI18185 bl<10> cbl<5> in1<78> in2<78> sl<10> vdd vss wl<78> / cell_PIM
XI18184 bl<10> cbl<5> in1<79> in2<79> sl<10> vdd vss wl<79> / cell_PIM
XI18838 bl<18> cbl<9> in1<123> in2<123> sl<18> vdd vss wl<123> / cell_PIM
XI18837 bl<18> cbl<9> in1<124> in2<124> sl<18> vdd vss wl<124> / cell_PIM
XI17533 bl<4> cbl<2> in1<65> in2<65> sl<4> vdd vss wl<65> / cell_PIM
XI17532 bl<4> cbl<2> in1<64> in2<64> sl<4> vdd vss wl<64> / cell_PIM
XI17531 bl<4> cbl<2> in1<63> in2<63> sl<4> vdd vss wl<63> / cell_PIM
XI18183 bl<10> cbl<5> in1<80> in2<80> sl<10> vdd vss wl<80> / cell_PIM
XI18182 bl<10> cbl<5> in1<81> in2<81> sl<10> vdd vss wl<81> / cell_PIM
XI18181 bl<10> cbl<5> in1<77> in2<77> sl<10> vdd vss wl<77> / cell_PIM
XI18831 bl<16> cbl<8> in1<127> in2<127> sl<16> vdd vss wl<127> / cell_PIM
XI18830 bl<16> cbl<8> in1<126> in2<126> sl<16> vdd vss wl<126> / cell_PIM
XI18829 bl<16> cbl<8> in1<125> in2<125> sl<16> vdd vss wl<125> / cell_PIM
XI18828 bl<16> cbl<8> in1<124> in2<124> sl<16> vdd vss wl<124> / cell_PIM
XI18827 bl<16> cbl<8> in1<123> in2<123> sl<16> vdd vss wl<123> / cell_PIM
XI18825 bl<14> cbl<7> in1<0> in2<0> sl<14> vdd vss wl<0> / cell_PIM
XI18175 bl<8> cbl<4> in1<81> in2<81> sl<8> vdd vss wl<81> / cell_PIM
XI18174 bl<8> cbl<4> in1<80> in2<80> sl<8> vdd vss wl<80> / cell_PIM
XI17526 bl<6> cbl<3> in1<69> in2<69> sl<6> vdd vss wl<69> / cell_PIM
XI17525 bl<6> cbl<3> in1<70> in2<70> sl<6> vdd vss wl<70> / cell_PIM
XI17524 bl<6> cbl<3> in1<71> in2<71> sl<6> vdd vss wl<71> / cell_PIM
XI17523 bl<6> cbl<3> in1<68> in2<68> sl<6> vdd vss wl<68> / cell_PIM
XI18173 bl<8> cbl<4> in1<79> in2<79> sl<8> vdd vss wl<79> / cell_PIM
XI18172 bl<8> cbl<4> in1<78> in2<78> sl<8> vdd vss wl<78> / cell_PIM
XI18171 bl<8> cbl<4> in1<77> in2<77> sl<8> vdd vss wl<77> / cell_PIM
XI18823 bl<12> cbl<6> in1<0> in2<0> sl<12> vdd vss wl<0> / cell_PIM
XI18821 bl<10> cbl<5> in1<0> in2<0> sl<10> vdd vss wl<0> / cell_PIM
XI18819 bl<8> cbl<4> in1<0> in2<0> sl<8> vdd vss wl<0> / cell_PIM
XI17518 bl<4> cbl<2> in1<71> in2<71> sl<4> vdd vss wl<71> / cell_PIM
XI17517 bl<4> cbl<2> in1<70> in2<70> sl<4> vdd vss wl<70> / cell_PIM
XI17516 bl<4> cbl<2> in1<69> in2<69> sl<4> vdd vss wl<69> / cell_PIM
XI17515 bl<4> cbl<2> in1<68> in2<68> sl<4> vdd vss wl<68> / cell_PIM
XI18165 bl<14> cbl<7> in1<83> in2<83> sl<14> vdd vss wl<83> / cell_PIM
XI18164 bl<14> cbl<7> in1<84> in2<84> sl<14> vdd vss wl<84> / cell_PIM
XI18814 bl<14> cbl<7> in1<1> in2<1> sl<14> vdd vss wl<1> / cell_PIM
XI17509 bl<6> cbl<3> in1<73> in2<73> sl<6> vdd vss wl<73> / cell_PIM
XI18163 bl<14> cbl<7> in1<85> in2<85> sl<14> vdd vss wl<85> / cell_PIM
XI18162 bl<14> cbl<7> in1<86> in2<86> sl<14> vdd vss wl<86> / cell_PIM
XI18161 bl<14> cbl<7> in1<82> in2<82> sl<14> vdd vss wl<82> / cell_PIM
XI18813 bl<14> cbl<7> in1<2> in2<2> sl<14> vdd vss wl<2> / cell_PIM
XI18812 bl<14> cbl<7> in1<3> in2<3> sl<14> vdd vss wl<3> / cell_PIM
XI18811 bl<14> cbl<7> in1<4> in2<4> sl<14> vdd vss wl<4> / cell_PIM
XI18806 bl<12> cbl<6> in1<4> in2<4> sl<12> vdd vss wl<4> / cell_PIM
XI18805 bl<12> cbl<6> in1<3> in2<3> sl<12> vdd vss wl<3> / cell_PIM
XI18804 bl<12> cbl<6> in1<2> in2<2> sl<12> vdd vss wl<2> / cell_PIM
XI18155 bl<12> cbl<6> in1<86> in2<86> sl<12> vdd vss wl<86> / cell_PIM
XI18154 bl<12> cbl<6> in1<85> in2<85> sl<12> vdd vss wl<85> / cell_PIM
XI17508 bl<6> cbl<3> in1<74> in2<74> sl<6> vdd vss wl<74> / cell_PIM
XI17507 bl<6> cbl<3> in1<75> in2<75> sl<6> vdd vss wl<75> / cell_PIM
XI17506 bl<6> cbl<3> in1<76> in2<76> sl<6> vdd vss wl<76> / cell_PIM
XI17505 bl<6> cbl<3> in1<72> in2<72> sl<6> vdd vss wl<72> / cell_PIM
XI17499 bl<4> cbl<2> in1<76> in2<76> sl<4> vdd vss wl<76> / cell_PIM
XI18153 bl<12> cbl<6> in1<84> in2<84> sl<12> vdd vss wl<84> / cell_PIM
XI18152 bl<12> cbl<6> in1<83> in2<83> sl<12> vdd vss wl<83> / cell_PIM
XI18151 bl<12> cbl<6> in1<82> in2<82> sl<12> vdd vss wl<82> / cell_PIM
XI18803 bl<12> cbl<6> in1<1> in2<1> sl<12> vdd vss wl<1> / cell_PIM
XI17498 bl<4> cbl<2> in1<75> in2<75> sl<4> vdd vss wl<75> / cell_PIM
XI17497 bl<4> cbl<2> in1<74> in2<74> sl<4> vdd vss wl<74> / cell_PIM
XI17496 bl<4> cbl<2> in1<73> in2<73> sl<4> vdd vss wl<73> / cell_PIM
XI17495 bl<4> cbl<2> in1<72> in2<72> sl<4> vdd vss wl<72> / cell_PIM
XI18145 bl<10> cbl<5> in1<83> in2<83> sl<10> vdd vss wl<83> / cell_PIM
XI18144 bl<10> cbl<5> in1<84> in2<84> sl<10> vdd vss wl<84> / cell_PIM
XI18798 bl<10> cbl<5> in1<1> in2<1> sl<10> vdd vss wl<1> / cell_PIM
XI18797 bl<10> cbl<5> in1<2> in2<2> sl<10> vdd vss wl<2> / cell_PIM
XI18796 bl<10> cbl<5> in1<3> in2<3> sl<10> vdd vss wl<3> / cell_PIM
XI18795 bl<10> cbl<5> in1<4> in2<4> sl<10> vdd vss wl<4> / cell_PIM
XI16906 bl<0> cbl<0> in1<127> in2<127> sl<0> vdd vss wl<127> / cell_PIM
XI16904 bl<0> cbl<0> in1<125> in2<125> sl<0> vdd vss wl<125> / cell_PIM
XI16903 bl<0> cbl<0> in1<124> in2<124> sl<0> vdd vss wl<124> / cell_PIM
XI16901 bl<0> cbl<0> in1<122> in2<122> sl<0> vdd vss wl<122> / cell_PIM
XI16900 bl<0> cbl<0> in1<121> in2<121> sl<0> vdd vss wl<121> / cell_PIM
XI16898 bl<0> cbl<0> in1<119> in2<119> sl<0> vdd vss wl<119> / cell_PIM
XI16897 bl<0> cbl<0> in1<118> in2<118> sl<0> vdd vss wl<118> / cell_PIM
XI16895 bl<0> cbl<0> in1<116> in2<116> sl<0> vdd vss wl<116> / cell_PIM
XI16894 bl<0> cbl<0> in1<115> in2<115> sl<0> vdd vss wl<115> / cell_PIM
XI16892 bl<0> cbl<0> in1<113> in2<113> sl<0> vdd vss wl<113> / cell_PIM
XI16891 bl<0> cbl<0> in1<112> in2<112> sl<0> vdd vss wl<112> / cell_PIM
XI16889 bl<0> cbl<0> in1<110> in2<110> sl<0> vdd vss wl<110> / cell_PIM
XI16888 bl<0> cbl<0> in1<109> in2<109> sl<0> vdd vss wl<109> / cell_PIM
XI16886 bl<0> cbl<0> in1<107> in2<107> sl<0> vdd vss wl<107> / cell_PIM
XI16885 bl<0> cbl<0> in1<106> in2<106> sl<0> vdd vss wl<106> / cell_PIM
XI16883 bl<0> cbl<0> in1<104> in2<104> sl<0> vdd vss wl<104> / cell_PIM
XI16882 bl<0> cbl<0> in1<103> in2<103> sl<0> vdd vss wl<103> / cell_PIM
XI16880 bl<0> cbl<0> in1<101> in2<101> sl<0> vdd vss wl<101> / cell_PIM
XI16879 bl<0> cbl<0> in1<100> in2<100> sl<0> vdd vss wl<100> / cell_PIM
XI16877 bl<0> cbl<0> in1<98> in2<98> sl<0> vdd vss wl<98> / cell_PIM
XI16876 bl<0> cbl<0> in1<97> in2<97> sl<0> vdd vss wl<97> / cell_PIM
XI25031 bl<60> cbl<30> vdd vdd sl<60> vdd vss vss / cell_PIM
XI25029 bl<58> cbl<29> vdd vdd sl<58> vdd vss vss / cell_PIM
XI25033 bl<62> cbl<31> vdd vdd sl<62> vdd vss vss / cell_PIM
XI25027 bl<56> cbl<28> vdd vdd sl<56> vdd vss vss / cell_PIM
XI25025 bl<54> cbl<27> vdd vdd sl<54> vdd vss vss / cell_PIM
XI24373 bl<58> cbl<29> in1<19> in2<19> sl<58> vdd vss wl<19> / cell_PIM
XI25021 bl<50> cbl<25> vdd vdd sl<50> vdd vss vss / cell_PIM
XI25019 bl<48> cbl<24> vdd vdd sl<48> vdd vss vss / cell_PIM
XI25023 bl<52> cbl<26> vdd vdd sl<52> vdd vss vss / cell_PIM
XI25017 bl<46> cbl<23> vdd vdd sl<46> vdd vss vss / cell_PIM
XI25015 bl<44> cbl<22> vdd vdd sl<44> vdd vss vss / cell_PIM
XI24363 bl<56> cbl<28> in1<20> in2<20> sl<56> vdd vss wl<20> / cell_PIM
XI25011 bl<40> cbl<20> vdd vdd sl<40> vdd vss vss / cell_PIM
XI25009 bl<38> cbl<19> vdd vdd sl<38> vdd vss vss / cell_PIM
XI25013 bl<42> cbl<21> vdd vdd sl<42> vdd vss vss / cell_PIM
XI25007 bl<36> cbl<18> vdd vdd sl<36> vdd vss vss / cell_PIM
XI25005 bl<34> cbl<17> vdd vdd sl<34> vdd vss vss / cell_PIM
XI24358 bl<54> cbl<27> in1<18> in2<18> sl<54> vdd vss wl<18> / cell_PIM
XI25001 bl<30> cbl<15> vdd vdd sl<30> vdd vss vss / cell_PIM
XI24999 bl<28> cbl<14> vdd vdd sl<28> vdd vss vss / cell_PIM
XI25003 bl<32> cbl<16> vdd vdd sl<32> vdd vss vss / cell_PIM
XI24348 bl<52> cbl<26> in1<21> in2<21> sl<52> vdd vss wl<21> / cell_PIM
XI24997 bl<26> cbl<13> vdd vdd sl<26> vdd vss vss / cell_PIM
XI24995 bl<24> cbl<12> vdd vdd sl<24> vdd vss vss / cell_PIM
XI24991 bl<20> cbl<10> vdd vdd sl<20> vdd vss vss / cell_PIM
XI24989 bl<18> cbl<9> vdd vdd sl<18> vdd vss vss / cell_PIM
XI24993 bl<22> cbl<11> vdd vdd sl<22> vdd vss vss / cell_PIM
XI24987 bl<16> cbl<8> vdd vdd sl<16> vdd vss vss / cell_PIM
XI24985 bl<14> cbl<7> vdd vdd sl<14> vdd vss vss / cell_PIM
XI24333 bl<48> cbl<24> in1<18> in2<18> sl<48> vdd vss wl<18> / cell_PIM
XI24981 bl<10> cbl<5> vdd vdd sl<10> vdd vss vss / cell_PIM
XI24979 bl<8> cbl<4> vdd vdd sl<8> vdd vss vss / cell_PIM
XI24983 bl<12> cbl<6> vdd vdd sl<12> vdd vss vss / cell_PIM
XI24977 bl<6> cbl<3> vdd vdd sl<6> vdd vss vss / cell_PIM
XI24975 bl<4> cbl<2> vdd vdd sl<4> vdd vss vss / cell_PIM
XI24323 bl<46> cbl<23> in1<20> in2<20> sl<46> vdd vss wl<20> / cell_PIM
XI24971 bl<0> cbl<0> vdd vdd sl<0> vdd vss vss / cell_PIM
XI24973 bl<2> cbl<1> vdd vdd sl<2> vdd vss vss / cell_PIM
XI24967 bl<62> cbl<31> in1<0> in2<0> sl<62> vdd vss wl<0> / cell_PIM
XI24966 bl<62> cbl<31> in1<1> in2<1> sl<62> vdd vss wl<1> / cell_PIM
XI24965 bl<62> cbl<31> in1<2> in2<2> sl<62> vdd vss wl<2> / cell_PIM
XI24318 bl<44> cbl<22> in1<19> in2<19> sl<44> vdd vss wl<19> / cell_PIM
XI24961 bl<60> cbl<30> in1<0> in2<0> sl<60> vdd vss wl<0> / cell_PIM
XI24960 bl<60> cbl<30> in1<2> in2<2> sl<60> vdd vss wl<2> / cell_PIM
XI24959 bl<60> cbl<30> in1<1> in2<1> sl<60> vdd vss wl<1> / cell_PIM
XI24308 bl<42> cbl<21> in1<21> in2<21> sl<42> vdd vss wl<21> / cell_PIM
XI24955 bl<58> cbl<29> in1<0> in2<0> sl<58> vdd vss wl<0> / cell_PIM
XI24954 bl<58> cbl<29> in1<1> in2<1> sl<58> vdd vss wl<1> / cell_PIM
XI24949 bl<56> cbl<28> in1<0> in2<0> sl<56> vdd vss wl<0> / cell_PIM
XI24953 bl<58> cbl<29> in1<2> in2<2> sl<58> vdd vss wl<2> / cell_PIM
XI24948 bl<56> cbl<28> in1<2> in2<2> sl<56> vdd vss wl<2> / cell_PIM
XI24947 bl<56> cbl<28> in1<1> in2<1> sl<56> vdd vss wl<1> / cell_PIM
XI24293 bl<38> cbl<19> in1<19> in2<19> sl<38> vdd vss wl<19> / cell_PIM
XI24942 bl<54> cbl<27> in1<1> in2<1> sl<54> vdd vss wl<1> / cell_PIM
XI24941 bl<54> cbl<27> in1<2> in2<2> sl<54> vdd vss wl<2> / cell_PIM
XI24943 bl<54> cbl<27> in1<0> in2<0> sl<54> vdd vss wl<0> / cell_PIM
XI24937 bl<52> cbl<26> in1<0> in2<0> sl<52> vdd vss wl<0> / cell_PIM
XI24936 bl<52> cbl<26> in1<2> in2<2> sl<52> vdd vss wl<2> / cell_PIM
XI24935 bl<52> cbl<26> in1<1> in2<1> sl<52> vdd vss wl<1> / cell_PIM
XI24283 bl<36> cbl<18> in1<20> in2<20> sl<36> vdd vss wl<20> / cell_PIM
XI24931 bl<50> cbl<25> in1<0> in2<0> sl<50> vdd vss wl<0> / cell_PIM
XI24930 bl<50> cbl<25> in1<1> in2<1> sl<50> vdd vss wl<1> / cell_PIM
XI24929 bl<50> cbl<25> in1<2> in2<2> sl<50> vdd vss wl<2> / cell_PIM
XI24925 bl<48> cbl<24> in1<0> in2<0> sl<48> vdd vss wl<0> / cell_PIM
XI24924 bl<48> cbl<24> in1<2> in2<2> sl<48> vdd vss wl<2> / cell_PIM
XI24278 bl<34> cbl<17> in1<18> in2<18> sl<34> vdd vss wl<18> / cell_PIM
XI24919 bl<46> cbl<23> in1<0> in2<0> sl<46> vdd vss wl<0> / cell_PIM
XI24923 bl<48> cbl<24> in1<1> in2<1> sl<48> vdd vss wl<1> / cell_PIM
XI24268 bl<32> cbl<16> in1<21> in2<21> sl<32> vdd vss wl<21> / cell_PIM
XI24917 bl<46> cbl<23> in1<2> in2<2> sl<46> vdd vss wl<2> / cell_PIM
XI24918 bl<46> cbl<23> in1<1> in2<1> sl<46> vdd vss wl<1> / cell_PIM
XI24912 bl<44> cbl<22> in1<2> in2<2> sl<44> vdd vss wl<2> / cell_PIM
XI24911 bl<44> cbl<22> in1<1> in2<1> sl<44> vdd vss wl<1> / cell_PIM
XI24913 bl<44> cbl<22> in1<0> in2<0> sl<44> vdd vss wl<0> / cell_PIM
XI24907 bl<42> cbl<21> in1<0> in2<0> sl<42> vdd vss wl<0> / cell_PIM
XI24906 bl<42> cbl<21> in1<1> in2<1> sl<42> vdd vss wl<1> / cell_PIM
XI24905 bl<42> cbl<21> in1<2> in2<2> sl<42> vdd vss wl<2> / cell_PIM
XI24258 bl<62> cbl<31> in1<26> in2<26> sl<62> vdd vss wl<26> / cell_PIM
XI24901 bl<40> cbl<20> in1<0> in2<0> sl<40> vdd vss wl<0> / cell_PIM
XI24900 bl<40> cbl<20> in1<2> in2<2> sl<40> vdd vss wl<2> / cell_PIM
XI24899 bl<40> cbl<20> in1<1> in2<1> sl<40> vdd vss wl<1> / cell_PIM
XI24248 bl<60> cbl<30> in1<26> in2<26> sl<60> vdd vss wl<26> / cell_PIM
XI24895 bl<38> cbl<19> in1<0> in2<0> sl<38> vdd vss wl<0> / cell_PIM
XI24894 bl<38> cbl<19> in1<1> in2<1> sl<38> vdd vss wl<1> / cell_PIM
XI24889 bl<36> cbl<18> in1<0> in2<0> sl<36> vdd vss wl<0> / cell_PIM
XI24893 bl<38> cbl<19> in1<2> in2<2> sl<38> vdd vss wl<2> / cell_PIM
XI24888 bl<36> cbl<18> in1<2> in2<2> sl<36> vdd vss wl<2> / cell_PIM
XI24887 bl<36> cbl<18> in1<1> in2<1> sl<36> vdd vss wl<1> / cell_PIM
XI24238 bl<58> cbl<29> in1<26> in2<26> sl<58> vdd vss wl<26> / cell_PIM
XI24882 bl<34> cbl<17> in1<1> in2<1> sl<34> vdd vss wl<1> / cell_PIM
XI24881 bl<34> cbl<17> in1<2> in2<2> sl<34> vdd vss wl<2> / cell_PIM
XI24883 bl<34> cbl<17> in1<0> in2<0> sl<34> vdd vss wl<0> / cell_PIM
XI24228 bl<56> cbl<28> in1<26> in2<26> sl<56> vdd vss wl<26> / cell_PIM
XI24877 bl<32> cbl<16> in1<0> in2<0> sl<32> vdd vss wl<0> / cell_PIM
XI24876 bl<32> cbl<16> in1<2> in2<2> sl<32> vdd vss wl<2> / cell_PIM
XI24875 bl<32> cbl<16> in1<1> in2<1> sl<32> vdd vss wl<1> / cell_PIM
XI22563 bl<62> cbl<31> in1<78> in2<78> sl<62> vdd vss wl<78> / cell_PIM
XI23733 bl<50> cbl<25> in1<38> in2<38> sl<50> vdd vss wl<38> / cell_PIM
XI23732 bl<50> cbl<25> in1<40> in2<40> sl<50> vdd vss wl<40> / cell_PIM
XI23731 bl<50> cbl<25> in1<39> in2<39> sl<50> vdd vss wl<39> / cell_PIM
XI24382 bl<60> cbl<30> in1<19> in2<19> sl<60> vdd vss wl<19> / cell_PIM
XI24381 bl<60> cbl<30> in1<18> in2<18> sl<60> vdd vss wl<18> / cell_PIM
XI24380 bl<60> cbl<30> in1<21> in2<21> sl<60> vdd vss wl<21> / cell_PIM
XI24379 bl<60> cbl<30> in1<20> in2<20> sl<60> vdd vss wl<20> / cell_PIM
XI24374 bl<58> cbl<29> in1<18> in2<18> sl<58> vdd vss wl<18> / cell_PIM
XI23726 bl<48> cbl<24> in1<38> in2<38> sl<48> vdd vss wl<38> / cell_PIM
XI23725 bl<48> cbl<24> in1<37> in2<37> sl<48> vdd vss wl<37> / cell_PIM
XI23724 bl<48> cbl<24> in1<40> in2<40> sl<48> vdd vss wl<40> / cell_PIM
XI23143 bl<56> cbl<28> in1<56> in2<56> sl<56> vdd vss wl<56> / cell_PIM
XI23142 bl<56> cbl<28> in1<57> in2<57> sl<56> vdd vss wl<57> / cell_PIM
XI23141 bl<56> cbl<28> in1<59> in2<59> sl<56> vdd vss wl<59> / cell_PIM
XI22553 bl<60> cbl<30> in1<79> in2<79> sl<60> vdd vss wl<79> / cell_PIM
XI23140 bl<56> cbl<28> in1<60> in2<60> sl<56> vdd vss wl<60> / cell_PIM
XI23139 bl<56> cbl<28> in1<58> in2<58> sl<56> vdd vss wl<58> / cell_PIM
XI23723 bl<48> cbl<24> in1<39> in2<39> sl<48> vdd vss wl<39> / cell_PIM
XI24372 bl<58> cbl<29> in1<21> in2<21> sl<58> vdd vss wl<21> / cell_PIM
XI24371 bl<58> cbl<29> in1<20> in2<20> sl<58> vdd vss wl<20> / cell_PIM
XI23133 bl<54> cbl<27> in1<56> in2<56> sl<54> vdd vss wl<56> / cell_PIM
XI23718 bl<46> cbl<23> in1<37> in2<37> sl<46> vdd vss wl<37> / cell_PIM
XI23717 bl<46> cbl<23> in1<38> in2<38> sl<46> vdd vss wl<38> / cell_PIM
XI23716 bl<46> cbl<23> in1<40> in2<40> sl<46> vdd vss wl<40> / cell_PIM
XI23715 bl<46> cbl<23> in1<39> in2<39> sl<46> vdd vss wl<39> / cell_PIM
XI24366 bl<56> cbl<28> in1<18> in2<18> sl<56> vdd vss wl<18> / cell_PIM
XI24365 bl<56> cbl<28> in1<19> in2<19> sl<56> vdd vss wl<19> / cell_PIM
XI24364 bl<56> cbl<28> in1<21> in2<21> sl<56> vdd vss wl<21> / cell_PIM
XI22543 bl<58> cbl<29> in1<78> in2<78> sl<58> vdd vss wl<78> / cell_PIM
XI23132 bl<54> cbl<27> in1<57> in2<57> sl<54> vdd vss wl<57> / cell_PIM
XI23131 bl<54> cbl<27> in1<59> in2<59> sl<54> vdd vss wl<59> / cell_PIM
XI23130 bl<54> cbl<27> in1<60> in2<60> sl<54> vdd vss wl<60> / cell_PIM
XI23129 bl<54> cbl<27> in1<58> in2<58> sl<54> vdd vss wl<58> / cell_PIM
XI23710 bl<44> cbl<22> in1<38> in2<38> sl<44> vdd vss wl<38> / cell_PIM
XI23709 bl<44> cbl<22> in1<37> in2<37> sl<44> vdd vss wl<37> / cell_PIM
XI24357 bl<54> cbl<27> in1<19> in2<19> sl<54> vdd vss wl<19> / cell_PIM
XI24356 bl<54> cbl<27> in1<21> in2<21> sl<54> vdd vss wl<21> / cell_PIM
XI24355 bl<54> cbl<27> in1<20> in2<20> sl<54> vdd vss wl<20> / cell_PIM
XI23708 bl<44> cbl<22> in1<40> in2<40> sl<44> vdd vss wl<40> / cell_PIM
XI23707 bl<44> cbl<22> in1<39> in2<39> sl<44> vdd vss wl<39> / cell_PIM
XI22533 bl<56> cbl<28> in1<78> in2<78> sl<56> vdd vss wl<78> / cell_PIM
XI23123 bl<52> cbl<26> in1<57> in2<57> sl<52> vdd vss wl<57> / cell_PIM
XI23122 bl<52> cbl<26> in1<56> in2<56> sl<52> vdd vss wl<56> / cell_PIM
XI23121 bl<52> cbl<26> in1<60> in2<60> sl<52> vdd vss wl<60> / cell_PIM
XI23702 bl<42> cbl<21> in1<37> in2<37> sl<42> vdd vss wl<37> / cell_PIM
XI23701 bl<42> cbl<21> in1<38> in2<38> sl<42> vdd vss wl<38> / cell_PIM
XI23700 bl<42> cbl<21> in1<40> in2<40> sl<42> vdd vss wl<40> / cell_PIM
XI23699 bl<42> cbl<21> in1<39> in2<39> sl<42> vdd vss wl<39> / cell_PIM
XI24350 bl<52> cbl<26> in1<19> in2<19> sl<52> vdd vss wl<19> / cell_PIM
XI24349 bl<52> cbl<26> in1<18> in2<18> sl<52> vdd vss wl<18> / cell_PIM
XI23120 bl<52> cbl<26> in1<59> in2<59> sl<52> vdd vss wl<59> / cell_PIM
XI23119 bl<52> cbl<26> in1<58> in2<58> sl<52> vdd vss wl<58> / cell_PIM
XI23694 bl<40> cbl<20> in1<37> in2<37> sl<40> vdd vss wl<37> / cell_PIM
XI24347 bl<52> cbl<26> in1<20> in2<20> sl<52> vdd vss wl<20> / cell_PIM
XI22523 bl<54> cbl<27> in1<78> in2<78> sl<54> vdd vss wl<78> / cell_PIM
XI23113 bl<50> cbl<25> in1<56> in2<56> sl<50> vdd vss wl<56> / cell_PIM
XI23693 bl<40> cbl<20> in1<38> in2<38> sl<40> vdd vss wl<38> / cell_PIM
XI23692 bl<40> cbl<20> in1<40> in2<40> sl<40> vdd vss wl<40> / cell_PIM
XI23691 bl<40> cbl<20> in1<39> in2<39> sl<40> vdd vss wl<39> / cell_PIM
XI24342 bl<50> cbl<25> in1<18> in2<18> sl<50> vdd vss wl<18> / cell_PIM
XI24341 bl<50> cbl<25> in1<19> in2<19> sl<50> vdd vss wl<19> / cell_PIM
XI24340 bl<50> cbl<25> in1<21> in2<21> sl<50> vdd vss wl<21> / cell_PIM
XI24339 bl<50> cbl<25> in1<20> in2<20> sl<50> vdd vss wl<20> / cell_PIM
XI24334 bl<48> cbl<24> in1<19> in2<19> sl<48> vdd vss wl<19> / cell_PIM
XI23686 bl<38> cbl<19> in1<37> in2<37> sl<38> vdd vss wl<37> / cell_PIM
XI23685 bl<38> cbl<19> in1<38> in2<38> sl<38> vdd vss wl<38> / cell_PIM
XI23684 bl<38> cbl<19> in1<40> in2<40> sl<38> vdd vss wl<40> / cell_PIM
XI23112 bl<50> cbl<25> in1<57> in2<57> sl<50> vdd vss wl<57> / cell_PIM
XI23111 bl<50> cbl<25> in1<59> in2<59> sl<50> vdd vss wl<59> / cell_PIM
XI23110 bl<50> cbl<25> in1<60> in2<60> sl<50> vdd vss wl<60> / cell_PIM
XI23109 bl<50> cbl<25> in1<58> in2<58> sl<50> vdd vss wl<58> / cell_PIM
XI22513 bl<52> cbl<26> in1<79> in2<79> sl<52> vdd vss wl<79> / cell_PIM
XI23683 bl<38> cbl<19> in1<39> in2<39> sl<38> vdd vss wl<39> / cell_PIM
XI24332 bl<48> cbl<24> in1<21> in2<21> sl<48> vdd vss wl<21> / cell_PIM
XI24331 bl<48> cbl<24> in1<20> in2<20> sl<48> vdd vss wl<20> / cell_PIM
XI23103 bl<48> cbl<24> in1<57> in2<57> sl<48> vdd vss wl<57> / cell_PIM
XI23102 bl<48> cbl<24> in1<56> in2<56> sl<48> vdd vss wl<56> / cell_PIM
XI23101 bl<48> cbl<24> in1<60> in2<60> sl<48> vdd vss wl<60> / cell_PIM
XI23678 bl<36> cbl<18> in1<38> in2<38> sl<36> vdd vss wl<38> / cell_PIM
XI23677 bl<36> cbl<18> in1<37> in2<37> sl<36> vdd vss wl<37> / cell_PIM
XI23676 bl<36> cbl<18> in1<40> in2<40> sl<36> vdd vss wl<40> / cell_PIM
XI23675 bl<36> cbl<18> in1<39> in2<39> sl<36> vdd vss wl<39> / cell_PIM
XI24326 bl<46> cbl<23> in1<18> in2<18> sl<46> vdd vss wl<18> / cell_PIM
XI24325 bl<46> cbl<23> in1<19> in2<19> sl<46> vdd vss wl<19> / cell_PIM
XI24324 bl<46> cbl<23> in1<21> in2<21> sl<46> vdd vss wl<21> / cell_PIM
XI22503 bl<50> cbl<25> in1<78> in2<78> sl<50> vdd vss wl<78> / cell_PIM
XI23100 bl<48> cbl<24> in1<59> in2<59> sl<48> vdd vss wl<59> / cell_PIM
XI23099 bl<48> cbl<24> in1<58> in2<58> sl<48> vdd vss wl<58> / cell_PIM
XI23670 bl<34> cbl<17> in1<37> in2<37> sl<34> vdd vss wl<37> / cell_PIM
XI23669 bl<34> cbl<17> in1<38> in2<38> sl<34> vdd vss wl<38> / cell_PIM
XI24317 bl<44> cbl<22> in1<18> in2<18> sl<44> vdd vss wl<18> / cell_PIM
XI24316 bl<44> cbl<22> in1<21> in2<21> sl<44> vdd vss wl<21> / cell_PIM
XI24315 bl<44> cbl<22> in1<20> in2<20> sl<44> vdd vss wl<20> / cell_PIM
XI23668 bl<34> cbl<17> in1<40> in2<40> sl<34> vdd vss wl<40> / cell_PIM
XI23667 bl<34> cbl<17> in1<39> in2<39> sl<34> vdd vss wl<39> / cell_PIM
XI23093 bl<46> cbl<23> in1<56> in2<56> sl<46> vdd vss wl<56> / cell_PIM
XI22493 bl<48> cbl<24> in1<79> in2<79> sl<48> vdd vss wl<79> / cell_PIM
XI23092 bl<46> cbl<23> in1<57> in2<57> sl<46> vdd vss wl<57> / cell_PIM
XI23091 bl<46> cbl<23> in1<59> in2<59> sl<46> vdd vss wl<59> / cell_PIM
XI23090 bl<46> cbl<23> in1<60> in2<60> sl<46> vdd vss wl<60> / cell_PIM
XI23089 bl<46> cbl<23> in1<58> in2<58> sl<46> vdd vss wl<58> / cell_PIM
XI23662 bl<32> cbl<16> in1<38> in2<38> sl<32> vdd vss wl<38> / cell_PIM
XI23661 bl<32> cbl<16> in1<37> in2<37> sl<32> vdd vss wl<37> / cell_PIM
XI23660 bl<32> cbl<16> in1<40> in2<40> sl<32> vdd vss wl<40> / cell_PIM
XI23659 bl<32> cbl<16> in1<39> in2<39> sl<32> vdd vss wl<39> / cell_PIM
XI24310 bl<42> cbl<21> in1<18> in2<18> sl<42> vdd vss wl<18> / cell_PIM
XI24309 bl<42> cbl<21> in1<19> in2<19> sl<42> vdd vss wl<19> / cell_PIM
XI24307 bl<42> cbl<21> in1<20> in2<20> sl<42> vdd vss wl<20> / cell_PIM
XI22483 bl<46> cbl<23> in1<78> in2<78> sl<46> vdd vss wl<78> / cell_PIM
XI23083 bl<44> cbl<22> in1<57> in2<57> sl<44> vdd vss wl<57> / cell_PIM
XI23082 bl<44> cbl<22> in1<56> in2<56> sl<44> vdd vss wl<56> / cell_PIM
XI23081 bl<44> cbl<22> in1<60> in2<60> sl<44> vdd vss wl<60> / cell_PIM
XI23653 bl<62> cbl<31> in1<41> in2<41> sl<62> vdd vss wl<41> / cell_PIM
XI23652 bl<62> cbl<31> in1<42> in2<42> sl<62> vdd vss wl<42> / cell_PIM
XI23651 bl<62> cbl<31> in1<43> in2<43> sl<62> vdd vss wl<43> / cell_PIM
XI23650 bl<62> cbl<31> in1<45> in2<45> sl<62> vdd vss wl<45> / cell_PIM
XI23649 bl<62> cbl<31> in1<44> in2<44> sl<62> vdd vss wl<44> / cell_PIM
XI24302 bl<40> cbl<20> in1<18> in2<18> sl<40> vdd vss wl<18> / cell_PIM
XI24301 bl<40> cbl<20> in1<19> in2<19> sl<40> vdd vss wl<19> / cell_PIM
XI24300 bl<40> cbl<20> in1<21> in2<21> sl<40> vdd vss wl<21> / cell_PIM
XI24299 bl<40> cbl<20> in1<20> in2<20> sl<40> vdd vss wl<20> / cell_PIM
XI24294 bl<38> cbl<19> in1<18> in2<18> sl<38> vdd vss wl<18> / cell_PIM
XI23080 bl<44> cbl<22> in1<59> in2<59> sl<44> vdd vss wl<59> / cell_PIM
XI23079 bl<44> cbl<22> in1<58> in2<58> sl<44> vdd vss wl<58> / cell_PIM
XI22473 bl<44> cbl<22> in1<79> in2<79> sl<44> vdd vss wl<79> / cell_PIM
XI23073 bl<42> cbl<21> in1<56> in2<56> sl<42> vdd vss wl<56> / cell_PIM
XI23643 bl<60> cbl<30> in1<43> in2<43> sl<60> vdd vss wl<43> / cell_PIM
XI23642 bl<60> cbl<30> in1<42> in2<42> sl<60> vdd vss wl<42> / cell_PIM
XI23641 bl<60> cbl<30> in1<41> in2<41> sl<60> vdd vss wl<41> / cell_PIM
XI23640 bl<60> cbl<30> in1<45> in2<45> sl<60> vdd vss wl<45> / cell_PIM
XI23639 bl<60> cbl<30> in1<44> in2<44> sl<60> vdd vss wl<44> / cell_PIM
XI24292 bl<38> cbl<19> in1<21> in2<21> sl<38> vdd vss wl<21> / cell_PIM
XI24291 bl<38> cbl<19> in1<20> in2<20> sl<38> vdd vss wl<20> / cell_PIM
XI23072 bl<42> cbl<21> in1<57> in2<57> sl<42> vdd vss wl<57> / cell_PIM
XI23071 bl<42> cbl<21> in1<59> in2<59> sl<42> vdd vss wl<59> / cell_PIM
XI23070 bl<42> cbl<21> in1<60> in2<60> sl<42> vdd vss wl<60> / cell_PIM
XI23069 bl<42> cbl<21> in1<58> in2<58> sl<42> vdd vss wl<58> / cell_PIM
XI24286 bl<36> cbl<18> in1<19> in2<19> sl<36> vdd vss wl<19> / cell_PIM
XI24285 bl<36> cbl<18> in1<18> in2<18> sl<36> vdd vss wl<18> / cell_PIM
XI24284 bl<36> cbl<18> in1<21> in2<21> sl<36> vdd vss wl<21> / cell_PIM
XI22463 bl<42> cbl<21> in1<78> in2<78> sl<42> vdd vss wl<78> / cell_PIM
XI23633 bl<58> cbl<29> in1<41> in2<41> sl<58> vdd vss wl<41> / cell_PIM
XI23632 bl<58> cbl<29> in1<42> in2<42> sl<58> vdd vss wl<42> / cell_PIM
XI23631 bl<58> cbl<29> in1<43> in2<43> sl<58> vdd vss wl<43> / cell_PIM
XI23630 bl<58> cbl<29> in1<45> in2<45> sl<58> vdd vss wl<45> / cell_PIM
XI23629 bl<58> cbl<29> in1<44> in2<44> sl<58> vdd vss wl<44> / cell_PIM
XI24277 bl<34> cbl<17> in1<19> in2<19> sl<34> vdd vss wl<19> / cell_PIM
XI24276 bl<34> cbl<17> in1<21> in2<21> sl<34> vdd vss wl<21> / cell_PIM
XI24275 bl<34> cbl<17> in1<20> in2<20> sl<34> vdd vss wl<20> / cell_PIM
XI23063 bl<40> cbl<20> in1<56> in2<56> sl<40> vdd vss wl<56> / cell_PIM
XI23062 bl<40> cbl<20> in1<57> in2<57> sl<40> vdd vss wl<57> / cell_PIM
XI23061 bl<40> cbl<20> in1<59> in2<59> sl<40> vdd vss wl<59> / cell_PIM
XI22453 bl<40> cbl<20> in1<78> in2<78> sl<40> vdd vss wl<78> / cell_PIM
XI23060 bl<40> cbl<20> in1<60> in2<60> sl<40> vdd vss wl<60> / cell_PIM
XI23059 bl<40> cbl<20> in1<58> in2<58> sl<40> vdd vss wl<58> / cell_PIM
XI23623 bl<56> cbl<28> in1<41> in2<41> sl<56> vdd vss wl<41> / cell_PIM
XI23622 bl<56> cbl<28> in1<42> in2<42> sl<56> vdd vss wl<42> / cell_PIM
XI23621 bl<56> cbl<28> in1<43> in2<43> sl<56> vdd vss wl<43> / cell_PIM
XI23620 bl<56> cbl<28> in1<45> in2<45> sl<56> vdd vss wl<45> / cell_PIM
XI23619 bl<56> cbl<28> in1<44> in2<44> sl<56> vdd vss wl<44> / cell_PIM
XI24270 bl<32> cbl<16> in1<19> in2<19> sl<32> vdd vss wl<19> / cell_PIM
XI24269 bl<32> cbl<16> in1<18> in2<18> sl<32> vdd vss wl<18> / cell_PIM
XI23053 bl<38> cbl<19> in1<56> in2<56> sl<38> vdd vss wl<56> / cell_PIM
XI24267 bl<32> cbl<16> in1<20> in2<20> sl<32> vdd vss wl<20> / cell_PIM
XI22443 bl<38> cbl<19> in1<78> in2<78> sl<38> vdd vss wl<78> / cell_PIM
XI23052 bl<38> cbl<19> in1<57> in2<57> sl<38> vdd vss wl<57> / cell_PIM
XI23051 bl<38> cbl<19> in1<59> in2<59> sl<38> vdd vss wl<59> / cell_PIM
XI23050 bl<38> cbl<19> in1<60> in2<60> sl<38> vdd vss wl<60> / cell_PIM
XI23049 bl<38> cbl<19> in1<58> in2<58> sl<38> vdd vss wl<58> / cell_PIM
XI23613 bl<54> cbl<27> in1<41> in2<41> sl<54> vdd vss wl<41> / cell_PIM
XI23612 bl<54> cbl<27> in1<42> in2<42> sl<54> vdd vss wl<42> / cell_PIM
XI23611 bl<54> cbl<27> in1<43> in2<43> sl<54> vdd vss wl<43> / cell_PIM
XI23610 bl<54> cbl<27> in1<45> in2<45> sl<54> vdd vss wl<45> / cell_PIM
XI23609 bl<54> cbl<27> in1<44> in2<44> sl<54> vdd vss wl<44> / cell_PIM
XI24261 bl<62> cbl<31> in1<22> in2<22> sl<62> vdd vss wl<22> / cell_PIM
XI24260 bl<62> cbl<31> in1<23> in2<23> sl<62> vdd vss wl<23> / cell_PIM
XI24259 bl<62> cbl<31> in1<24> in2<24> sl<62> vdd vss wl<24> / cell_PIM
XI24257 bl<62> cbl<31> in1<25> in2<25> sl<62> vdd vss wl<25> / cell_PIM
XI22433 bl<36> cbl<18> in1<79> in2<79> sl<36> vdd vss wl<79> / cell_PIM
XI23043 bl<36> cbl<18> in1<57> in2<57> sl<36> vdd vss wl<57> / cell_PIM
XI23042 bl<36> cbl<18> in1<56> in2<56> sl<36> vdd vss wl<56> / cell_PIM
XI23041 bl<36> cbl<18> in1<60> in2<60> sl<36> vdd vss wl<60> / cell_PIM
XI23603 bl<52> cbl<26> in1<43> in2<43> sl<52> vdd vss wl<43> / cell_PIM
XI23602 bl<52> cbl<26> in1<42> in2<42> sl<52> vdd vss wl<42> / cell_PIM
XI23601 bl<52> cbl<26> in1<41> in2<41> sl<52> vdd vss wl<41> / cell_PIM
XI23600 bl<52> cbl<26> in1<45> in2<45> sl<52> vdd vss wl<45> / cell_PIM
XI23599 bl<52> cbl<26> in1<44> in2<44> sl<52> vdd vss wl<44> / cell_PIM
XI24251 bl<60> cbl<30> in1<24> in2<24> sl<60> vdd vss wl<24> / cell_PIM
XI24250 bl<60> cbl<30> in1<23> in2<23> sl<60> vdd vss wl<23> / cell_PIM
XI24249 bl<60> cbl<30> in1<22> in2<22> sl<60> vdd vss wl<22> / cell_PIM
XI23040 bl<36> cbl<18> in1<59> in2<59> sl<36> vdd vss wl<59> / cell_PIM
XI23039 bl<36> cbl<18> in1<58> in2<58> sl<36> vdd vss wl<58> / cell_PIM
XI24247 bl<60> cbl<30> in1<25> in2<25> sl<60> vdd vss wl<25> / cell_PIM
XI22423 bl<34> cbl<17> in1<78> in2<78> sl<34> vdd vss wl<78> / cell_PIM
XI23033 bl<34> cbl<17> in1<56> in2<56> sl<34> vdd vss wl<56> / cell_PIM
XI23593 bl<50> cbl<25> in1<41> in2<41> sl<50> vdd vss wl<41> / cell_PIM
XI23592 bl<50> cbl<25> in1<42> in2<42> sl<50> vdd vss wl<42> / cell_PIM
XI23591 bl<50> cbl<25> in1<43> in2<43> sl<50> vdd vss wl<43> / cell_PIM
XI23590 bl<50> cbl<25> in1<45> in2<45> sl<50> vdd vss wl<45> / cell_PIM
XI23589 bl<50> cbl<25> in1<44> in2<44> sl<50> vdd vss wl<44> / cell_PIM
XI24241 bl<58> cbl<29> in1<22> in2<22> sl<58> vdd vss wl<22> / cell_PIM
XI24240 bl<58> cbl<29> in1<23> in2<23> sl<58> vdd vss wl<23> / cell_PIM
XI24239 bl<58> cbl<29> in1<24> in2<24> sl<58> vdd vss wl<24> / cell_PIM
XI24237 bl<58> cbl<29> in1<25> in2<25> sl<58> vdd vss wl<25> / cell_PIM
XI23032 bl<34> cbl<17> in1<57> in2<57> sl<34> vdd vss wl<57> / cell_PIM
XI23031 bl<34> cbl<17> in1<59> in2<59> sl<34> vdd vss wl<59> / cell_PIM
XI23030 bl<34> cbl<17> in1<60> in2<60> sl<34> vdd vss wl<60> / cell_PIM
XI23029 bl<34> cbl<17> in1<58> in2<58> sl<34> vdd vss wl<58> / cell_PIM
XI22413 bl<32> cbl<16> in1<79> in2<79> sl<32> vdd vss wl<79> / cell_PIM
XI23583 bl<48> cbl<24> in1<43> in2<43> sl<48> vdd vss wl<43> / cell_PIM
XI23582 bl<48> cbl<24> in1<42> in2<42> sl<48> vdd vss wl<42> / cell_PIM
XI23581 bl<48> cbl<24> in1<41> in2<41> sl<48> vdd vss wl<41> / cell_PIM
XI23580 bl<48> cbl<24> in1<45> in2<45> sl<48> vdd vss wl<45> / cell_PIM
XI23579 bl<48> cbl<24> in1<44> in2<44> sl<48> vdd vss wl<44> / cell_PIM
XI24231 bl<56> cbl<28> in1<22> in2<22> sl<56> vdd vss wl<22> / cell_PIM
XI24230 bl<56> cbl<28> in1<23> in2<23> sl<56> vdd vss wl<23> / cell_PIM
XI24229 bl<56> cbl<28> in1<24> in2<24> sl<56> vdd vss wl<24> / cell_PIM
XI23023 bl<32> cbl<16> in1<57> in2<57> sl<32> vdd vss wl<57> / cell_PIM
XI23022 bl<32> cbl<16> in1<56> in2<56> sl<32> vdd vss wl<56> / cell_PIM
XI23021 bl<32> cbl<16> in1<60> in2<60> sl<32> vdd vss wl<60> / cell_PIM
XI24227 bl<56> cbl<28> in1<25> in2<25> sl<56> vdd vss wl<25> / cell_PIM
XI21259 bl<44> cbl<22> in1<115> in2<115> sl<44> vdd vss wl<115> / cell_PIM
XI21913 bl<54> cbl<27> in1<96> in2<96> sl<54> vdd vss wl<96> / cell_PIM
XI22562 bl<62> cbl<31> in1<79> in2<79> sl<62> vdd vss wl<79> / cell_PIM
XI22561 bl<62> cbl<31> in1<77> in2<77> sl<62> vdd vss wl<77> / cell_PIM
XI22555 bl<60> cbl<30> in1<76> in2<76> sl<60> vdd vss wl<76> / cell_PIM
XI21907 bl<52> cbl<26> in1<95> in2<95> sl<52> vdd vss wl<95> / cell_PIM
XI21906 bl<52> cbl<26> in1<94> in2<94> sl<52> vdd vss wl<94> / cell_PIM
XI21905 bl<52> cbl<26> in1<98> in2<98> sl<52> vdd vss wl<98> / cell_PIM
XI21904 bl<52> cbl<26> in1<97> in2<97> sl<52> vdd vss wl<97> / cell_PIM
XI21258 bl<44> cbl<22> in1<114> in2<114> sl<44> vdd vss wl<114> / cell_PIM
XI21257 bl<44> cbl<22> in1<113> in2<113> sl<44> vdd vss wl<113> / cell_PIM
XI21256 bl<44> cbl<22> in1<117> in2<117> sl<44> vdd vss wl<117> / cell_PIM
XI21255 bl<44> cbl<22> in1<116> in2<116> sl<44> vdd vss wl<116> / cell_PIM
XI22554 bl<60> cbl<30> in1<75> in2<75> sl<60> vdd vss wl<75> / cell_PIM
XI21249 bl<42> cbl<21> in1<113> in2<113> sl<42> vdd vss wl<113> / cell_PIM
XI21903 bl<52> cbl<26> in1<96> in2<96> sl<52> vdd vss wl<96> / cell_PIM
XI22552 bl<60> cbl<30> in1<78> in2<78> sl<60> vdd vss wl<78> / cell_PIM
XI22551 bl<60> cbl<30> in1<77> in2<77> sl<60> vdd vss wl<77> / cell_PIM
XI21248 bl<42> cbl<21> in1<114> in2<114> sl<42> vdd vss wl<114> / cell_PIM
XI21247 bl<42> cbl<21> in1<115> in2<115> sl<42> vdd vss wl<115> / cell_PIM
XI21246 bl<42> cbl<21> in1<117> in2<117> sl<42> vdd vss wl<117> / cell_PIM
XI21245 bl<42> cbl<21> in1<116> in2<116> sl<42> vdd vss wl<116> / cell_PIM
XI21897 bl<50> cbl<25> in1<94> in2<94> sl<50> vdd vss wl<94> / cell_PIM
XI21896 bl<50> cbl<25> in1<95> in2<95> sl<50> vdd vss wl<95> / cell_PIM
XI21895 bl<50> cbl<25> in1<97> in2<97> sl<50> vdd vss wl<97> / cell_PIM
XI21894 bl<50> cbl<25> in1<98> in2<98> sl<50> vdd vss wl<98> / cell_PIM
XI22545 bl<58> cbl<29> in1<75> in2<75> sl<58> vdd vss wl<75> / cell_PIM
XI22544 bl<58> cbl<29> in1<76> in2<76> sl<58> vdd vss wl<76> / cell_PIM
XI21239 bl<40> cbl<20> in1<113> in2<113> sl<40> vdd vss wl<113> / cell_PIM
XI21893 bl<50> cbl<25> in1<96> in2<96> sl<50> vdd vss wl<96> / cell_PIM
XI22542 bl<58> cbl<29> in1<79> in2<79> sl<58> vdd vss wl<79> / cell_PIM
XI22541 bl<58> cbl<29> in1<77> in2<77> sl<58> vdd vss wl<77> / cell_PIM
XI22535 bl<56> cbl<28> in1<75> in2<75> sl<56> vdd vss wl<75> / cell_PIM
XI21887 bl<48> cbl<24> in1<95> in2<95> sl<48> vdd vss wl<95> / cell_PIM
XI21886 bl<48> cbl<24> in1<94> in2<94> sl<48> vdd vss wl<94> / cell_PIM
XI21885 bl<48> cbl<24> in1<98> in2<98> sl<48> vdd vss wl<98> / cell_PIM
XI21884 bl<48> cbl<24> in1<97> in2<97> sl<48> vdd vss wl<97> / cell_PIM
XI21238 bl<40> cbl<20> in1<114> in2<114> sl<40> vdd vss wl<114> / cell_PIM
XI21237 bl<40> cbl<20> in1<115> in2<115> sl<40> vdd vss wl<115> / cell_PIM
XI21236 bl<40> cbl<20> in1<117> in2<117> sl<40> vdd vss wl<117> / cell_PIM
XI21235 bl<40> cbl<20> in1<116> in2<116> sl<40> vdd vss wl<116> / cell_PIM
XI22534 bl<56> cbl<28> in1<76> in2<76> sl<56> vdd vss wl<76> / cell_PIM
XI21229 bl<38> cbl<19> in1<113> in2<113> sl<38> vdd vss wl<113> / cell_PIM
XI21883 bl<48> cbl<24> in1<96> in2<96> sl<48> vdd vss wl<96> / cell_PIM
XI22532 bl<56> cbl<28> in1<79> in2<79> sl<56> vdd vss wl<79> / cell_PIM
XI22531 bl<56> cbl<28> in1<77> in2<77> sl<56> vdd vss wl<77> / cell_PIM
XI21228 bl<38> cbl<19> in1<114> in2<114> sl<38> vdd vss wl<114> / cell_PIM
XI21227 bl<38> cbl<19> in1<115> in2<115> sl<38> vdd vss wl<115> / cell_PIM
XI21226 bl<38> cbl<19> in1<117> in2<117> sl<38> vdd vss wl<117> / cell_PIM
XI21225 bl<38> cbl<19> in1<116> in2<116> sl<38> vdd vss wl<116> / cell_PIM
XI21877 bl<46> cbl<23> in1<94> in2<94> sl<46> vdd vss wl<94> / cell_PIM
XI21876 bl<46> cbl<23> in1<95> in2<95> sl<46> vdd vss wl<95> / cell_PIM
XI21875 bl<46> cbl<23> in1<97> in2<97> sl<46> vdd vss wl<97> / cell_PIM
XI21874 bl<46> cbl<23> in1<98> in2<98> sl<46> vdd vss wl<98> / cell_PIM
XI22525 bl<54> cbl<27> in1<75> in2<75> sl<54> vdd vss wl<75> / cell_PIM
XI22524 bl<54> cbl<27> in1<76> in2<76> sl<54> vdd vss wl<76> / cell_PIM
XI21219 bl<36> cbl<18> in1<115> in2<115> sl<36> vdd vss wl<115> / cell_PIM
XI21873 bl<46> cbl<23> in1<96> in2<96> sl<46> vdd vss wl<96> / cell_PIM
XI22522 bl<54> cbl<27> in1<79> in2<79> sl<54> vdd vss wl<79> / cell_PIM
XI22521 bl<54> cbl<27> in1<77> in2<77> sl<54> vdd vss wl<77> / cell_PIM
XI22515 bl<52> cbl<26> in1<76> in2<76> sl<52> vdd vss wl<76> / cell_PIM
XI21867 bl<44> cbl<22> in1<95> in2<95> sl<44> vdd vss wl<95> / cell_PIM
XI21866 bl<44> cbl<22> in1<94> in2<94> sl<44> vdd vss wl<94> / cell_PIM
XI21865 bl<44> cbl<22> in1<98> in2<98> sl<44> vdd vss wl<98> / cell_PIM
XI21864 bl<44> cbl<22> in1<97> in2<97> sl<44> vdd vss wl<97> / cell_PIM
XI21218 bl<36> cbl<18> in1<114> in2<114> sl<36> vdd vss wl<114> / cell_PIM
XI21217 bl<36> cbl<18> in1<113> in2<113> sl<36> vdd vss wl<113> / cell_PIM
XI21216 bl<36> cbl<18> in1<117> in2<117> sl<36> vdd vss wl<117> / cell_PIM
XI21215 bl<36> cbl<18> in1<116> in2<116> sl<36> vdd vss wl<116> / cell_PIM
XI22514 bl<52> cbl<26> in1<75> in2<75> sl<52> vdd vss wl<75> / cell_PIM
XI21209 bl<34> cbl<17> in1<113> in2<113> sl<34> vdd vss wl<113> / cell_PIM
XI21863 bl<44> cbl<22> in1<96> in2<96> sl<44> vdd vss wl<96> / cell_PIM
XI22512 bl<52> cbl<26> in1<78> in2<78> sl<52> vdd vss wl<78> / cell_PIM
XI22511 bl<52> cbl<26> in1<77> in2<77> sl<52> vdd vss wl<77> / cell_PIM
XI21208 bl<34> cbl<17> in1<114> in2<114> sl<34> vdd vss wl<114> / cell_PIM
XI21207 bl<34> cbl<17> in1<115> in2<115> sl<34> vdd vss wl<115> / cell_PIM
XI21206 bl<34> cbl<17> in1<117> in2<117> sl<34> vdd vss wl<117> / cell_PIM
XI21205 bl<34> cbl<17> in1<116> in2<116> sl<34> vdd vss wl<116> / cell_PIM
XI21857 bl<42> cbl<21> in1<94> in2<94> sl<42> vdd vss wl<94> / cell_PIM
XI21856 bl<42> cbl<21> in1<95> in2<95> sl<42> vdd vss wl<95> / cell_PIM
XI21855 bl<42> cbl<21> in1<97> in2<97> sl<42> vdd vss wl<97> / cell_PIM
XI21854 bl<42> cbl<21> in1<98> in2<98> sl<42> vdd vss wl<98> / cell_PIM
XI22505 bl<50> cbl<25> in1<75> in2<75> sl<50> vdd vss wl<75> / cell_PIM
XI22504 bl<50> cbl<25> in1<76> in2<76> sl<50> vdd vss wl<76> / cell_PIM
XI21199 bl<32> cbl<16> in1<115> in2<115> sl<32> vdd vss wl<115> / cell_PIM
XI21853 bl<42> cbl<21> in1<96> in2<96> sl<42> vdd vss wl<96> / cell_PIM
XI22502 bl<50> cbl<25> in1<79> in2<79> sl<50> vdd vss wl<79> / cell_PIM
XI22501 bl<50> cbl<25> in1<77> in2<77> sl<50> vdd vss wl<77> / cell_PIM
XI22495 bl<48> cbl<24> in1<76> in2<76> sl<48> vdd vss wl<76> / cell_PIM
XI21847 bl<40> cbl<20> in1<94> in2<94> sl<40> vdd vss wl<94> / cell_PIM
XI21846 bl<40> cbl<20> in1<95> in2<95> sl<40> vdd vss wl<95> / cell_PIM
XI21845 bl<40> cbl<20> in1<97> in2<97> sl<40> vdd vss wl<97> / cell_PIM
XI21844 bl<40> cbl<20> in1<98> in2<98> sl<40> vdd vss wl<98> / cell_PIM
XI21198 bl<32> cbl<16> in1<114> in2<114> sl<32> vdd vss wl<114> / cell_PIM
XI21197 bl<32> cbl<16> in1<113> in2<113> sl<32> vdd vss wl<113> / cell_PIM
XI21196 bl<32> cbl<16> in1<117> in2<117> sl<32> vdd vss wl<117> / cell_PIM
XI21195 bl<32> cbl<16> in1<116> in2<116> sl<32> vdd vss wl<116> / cell_PIM
XI22494 bl<48> cbl<24> in1<75> in2<75> sl<48> vdd vss wl<75> / cell_PIM
XI21189 bl<62> cbl<31> in1<118> in2<118> sl<62> vdd vss wl<118> / cell_PIM
XI21843 bl<40> cbl<20> in1<96> in2<96> sl<40> vdd vss wl<96> / cell_PIM
XI22492 bl<48> cbl<24> in1<78> in2<78> sl<48> vdd vss wl<78> / cell_PIM
XI22491 bl<48> cbl<24> in1<77> in2<77> sl<48> vdd vss wl<77> / cell_PIM
XI21188 bl<62> cbl<31> in1<119> in2<119> sl<62> vdd vss wl<119> / cell_PIM
XI21187 bl<62> cbl<31> in1<121> in2<121> sl<62> vdd vss wl<121> / cell_PIM
XI21186 bl<62> cbl<31> in1<122> in2<122> sl<62> vdd vss wl<122> / cell_PIM
XI21185 bl<62> cbl<31> in1<120> in2<120> sl<62> vdd vss wl<120> / cell_PIM
XI21837 bl<38> cbl<19> in1<94> in2<94> sl<38> vdd vss wl<94> / cell_PIM
XI21836 bl<38> cbl<19> in1<95> in2<95> sl<38> vdd vss wl<95> / cell_PIM
XI21835 bl<38> cbl<19> in1<97> in2<97> sl<38> vdd vss wl<97> / cell_PIM
XI21834 bl<38> cbl<19> in1<98> in2<98> sl<38> vdd vss wl<98> / cell_PIM
XI22485 bl<46> cbl<23> in1<75> in2<75> sl<46> vdd vss wl<75> / cell_PIM
XI22484 bl<46> cbl<23> in1<76> in2<76> sl<46> vdd vss wl<76> / cell_PIM
XI21179 bl<60> cbl<30> in1<119> in2<119> sl<60> vdd vss wl<119> / cell_PIM
XI21833 bl<38> cbl<19> in1<96> in2<96> sl<38> vdd vss wl<96> / cell_PIM
XI22482 bl<46> cbl<23> in1<79> in2<79> sl<46> vdd vss wl<79> / cell_PIM
XI22481 bl<46> cbl<23> in1<77> in2<77> sl<46> vdd vss wl<77> / cell_PIM
XI22475 bl<44> cbl<22> in1<76> in2<76> sl<44> vdd vss wl<76> / cell_PIM
XI21827 bl<36> cbl<18> in1<95> in2<95> sl<36> vdd vss wl<95> / cell_PIM
XI21826 bl<36> cbl<18> in1<94> in2<94> sl<36> vdd vss wl<94> / cell_PIM
XI21825 bl<36> cbl<18> in1<98> in2<98> sl<36> vdd vss wl<98> / cell_PIM
XI21824 bl<36> cbl<18> in1<97> in2<97> sl<36> vdd vss wl<97> / cell_PIM
XI21178 bl<60> cbl<30> in1<118> in2<118> sl<60> vdd vss wl<118> / cell_PIM
XI21177 bl<60> cbl<30> in1<122> in2<122> sl<60> vdd vss wl<122> / cell_PIM
XI21176 bl<60> cbl<30> in1<121> in2<121> sl<60> vdd vss wl<121> / cell_PIM
XI21175 bl<60> cbl<30> in1<120> in2<120> sl<60> vdd vss wl<120> / cell_PIM
XI22474 bl<44> cbl<22> in1<75> in2<75> sl<44> vdd vss wl<75> / cell_PIM
XI21169 bl<58> cbl<29> in1<118> in2<118> sl<58> vdd vss wl<118> / cell_PIM
XI21823 bl<36> cbl<18> in1<96> in2<96> sl<36> vdd vss wl<96> / cell_PIM
XI22472 bl<44> cbl<22> in1<78> in2<78> sl<44> vdd vss wl<78> / cell_PIM
XI22471 bl<44> cbl<22> in1<77> in2<77> sl<44> vdd vss wl<77> / cell_PIM
XI21168 bl<58> cbl<29> in1<119> in2<119> sl<58> vdd vss wl<119> / cell_PIM
XI21167 bl<58> cbl<29> in1<121> in2<121> sl<58> vdd vss wl<121> / cell_PIM
XI21166 bl<58> cbl<29> in1<122> in2<122> sl<58> vdd vss wl<122> / cell_PIM
XI21165 bl<58> cbl<29> in1<120> in2<120> sl<58> vdd vss wl<120> / cell_PIM
XI21817 bl<34> cbl<17> in1<94> in2<94> sl<34> vdd vss wl<94> / cell_PIM
XI21816 bl<34> cbl<17> in1<95> in2<95> sl<34> vdd vss wl<95> / cell_PIM
XI21815 bl<34> cbl<17> in1<97> in2<97> sl<34> vdd vss wl<97> / cell_PIM
XI21814 bl<34> cbl<17> in1<98> in2<98> sl<34> vdd vss wl<98> / cell_PIM
XI22465 bl<42> cbl<21> in1<75> in2<75> sl<42> vdd vss wl<75> / cell_PIM
XI22464 bl<42> cbl<21> in1<76> in2<76> sl<42> vdd vss wl<76> / cell_PIM
XI21159 bl<56> cbl<28> in1<118> in2<118> sl<56> vdd vss wl<118> / cell_PIM
XI21813 bl<34> cbl<17> in1<96> in2<96> sl<34> vdd vss wl<96> / cell_PIM
XI22462 bl<42> cbl<21> in1<79> in2<79> sl<42> vdd vss wl<79> / cell_PIM
XI22461 bl<42> cbl<21> in1<77> in2<77> sl<42> vdd vss wl<77> / cell_PIM
XI22455 bl<40> cbl<20> in1<75> in2<75> sl<40> vdd vss wl<75> / cell_PIM
XI21807 bl<32> cbl<16> in1<95> in2<95> sl<32> vdd vss wl<95> / cell_PIM
XI21806 bl<32> cbl<16> in1<94> in2<94> sl<32> vdd vss wl<94> / cell_PIM
XI21805 bl<32> cbl<16> in1<98> in2<98> sl<32> vdd vss wl<98> / cell_PIM
XI21804 bl<32> cbl<16> in1<97> in2<97> sl<32> vdd vss wl<97> / cell_PIM
XI21158 bl<56> cbl<28> in1<119> in2<119> sl<56> vdd vss wl<119> / cell_PIM
XI21157 bl<56> cbl<28> in1<121> in2<121> sl<56> vdd vss wl<121> / cell_PIM
XI21156 bl<56> cbl<28> in1<122> in2<122> sl<56> vdd vss wl<122> / cell_PIM
XI21155 bl<56> cbl<28> in1<120> in2<120> sl<56> vdd vss wl<120> / cell_PIM
XI22454 bl<40> cbl<20> in1<76> in2<76> sl<40> vdd vss wl<76> / cell_PIM
XI21149 bl<54> cbl<27> in1<118> in2<118> sl<54> vdd vss wl<118> / cell_PIM
XI21803 bl<32> cbl<16> in1<96> in2<96> sl<32> vdd vss wl<96> / cell_PIM
XI22452 bl<40> cbl<20> in1<79> in2<79> sl<40> vdd vss wl<79> / cell_PIM
XI22451 bl<40> cbl<20> in1<77> in2<77> sl<40> vdd vss wl<77> / cell_PIM
XI21148 bl<54> cbl<27> in1<119> in2<119> sl<54> vdd vss wl<119> / cell_PIM
XI21147 bl<54> cbl<27> in1<121> in2<121> sl<54> vdd vss wl<121> / cell_PIM
XI21146 bl<54> cbl<27> in1<122> in2<122> sl<54> vdd vss wl<122> / cell_PIM
XI21145 bl<54> cbl<27> in1<120> in2<120> sl<54> vdd vss wl<120> / cell_PIM
XI21797 bl<62> cbl<31> in1<99> in2<99> sl<62> vdd vss wl<99> / cell_PIM
XI21796 bl<62> cbl<31> in1<100> in2<100> sl<62> vdd vss wl<100> / cell_PIM
XI21795 bl<62> cbl<31> in1<102> in2<102> sl<62> vdd vss wl<102> / cell_PIM
XI21794 bl<62> cbl<31> in1<103> in2<103> sl<62> vdd vss wl<103> / cell_PIM
XI22445 bl<38> cbl<19> in1<75> in2<75> sl<38> vdd vss wl<75> / cell_PIM
XI22444 bl<38> cbl<19> in1<76> in2<76> sl<38> vdd vss wl<76> / cell_PIM
XI21139 bl<52> cbl<26> in1<119> in2<119> sl<52> vdd vss wl<119> / cell_PIM
XI21793 bl<62> cbl<31> in1<101> in2<101> sl<62> vdd vss wl<101> / cell_PIM
XI22442 bl<38> cbl<19> in1<79> in2<79> sl<38> vdd vss wl<79> / cell_PIM
XI22441 bl<38> cbl<19> in1<77> in2<77> sl<38> vdd vss wl<77> / cell_PIM
XI22435 bl<36> cbl<18> in1<76> in2<76> sl<36> vdd vss wl<76> / cell_PIM
XI21787 bl<60> cbl<30> in1<100> in2<100> sl<60> vdd vss wl<100> / cell_PIM
XI21786 bl<60> cbl<30> in1<99> in2<99> sl<60> vdd vss wl<99> / cell_PIM
XI21785 bl<60> cbl<30> in1<103> in2<103> sl<60> vdd vss wl<103> / cell_PIM
XI21784 bl<60> cbl<30> in1<102> in2<102> sl<60> vdd vss wl<102> / cell_PIM
XI21138 bl<52> cbl<26> in1<118> in2<118> sl<52> vdd vss wl<118> / cell_PIM
XI21137 bl<52> cbl<26> in1<122> in2<122> sl<52> vdd vss wl<122> / cell_PIM
XI21136 bl<52> cbl<26> in1<121> in2<121> sl<52> vdd vss wl<121> / cell_PIM
XI21135 bl<52> cbl<26> in1<120> in2<120> sl<52> vdd vss wl<120> / cell_PIM
XI22434 bl<36> cbl<18> in1<75> in2<75> sl<36> vdd vss wl<75> / cell_PIM
XI21129 bl<50> cbl<25> in1<118> in2<118> sl<50> vdd vss wl<118> / cell_PIM
XI21783 bl<60> cbl<30> in1<101> in2<101> sl<60> vdd vss wl<101> / cell_PIM
XI22432 bl<36> cbl<18> in1<78> in2<78> sl<36> vdd vss wl<78> / cell_PIM
XI22431 bl<36> cbl<18> in1<77> in2<77> sl<36> vdd vss wl<77> / cell_PIM
XI21128 bl<50> cbl<25> in1<119> in2<119> sl<50> vdd vss wl<119> / cell_PIM
XI21127 bl<50> cbl<25> in1<121> in2<121> sl<50> vdd vss wl<121> / cell_PIM
XI21126 bl<50> cbl<25> in1<122> in2<122> sl<50> vdd vss wl<122> / cell_PIM
XI21125 bl<50> cbl<25> in1<120> in2<120> sl<50> vdd vss wl<120> / cell_PIM
XI21777 bl<58> cbl<29> in1<99> in2<99> sl<58> vdd vss wl<99> / cell_PIM
XI21776 bl<58> cbl<29> in1<100> in2<100> sl<58> vdd vss wl<100> / cell_PIM
XI21775 bl<58> cbl<29> in1<102> in2<102> sl<58> vdd vss wl<102> / cell_PIM
XI21774 bl<58> cbl<29> in1<103> in2<103> sl<58> vdd vss wl<103> / cell_PIM
XI22425 bl<34> cbl<17> in1<75> in2<75> sl<34> vdd vss wl<75> / cell_PIM
XI22424 bl<34> cbl<17> in1<76> in2<76> sl<34> vdd vss wl<76> / cell_PIM
XI21119 bl<48> cbl<24> in1<119> in2<119> sl<48> vdd vss wl<119> / cell_PIM
XI21773 bl<58> cbl<29> in1<101> in2<101> sl<58> vdd vss wl<101> / cell_PIM
XI22422 bl<34> cbl<17> in1<79> in2<79> sl<34> vdd vss wl<79> / cell_PIM
XI22421 bl<34> cbl<17> in1<77> in2<77> sl<34> vdd vss wl<77> / cell_PIM
XI22415 bl<32> cbl<16> in1<76> in2<76> sl<32> vdd vss wl<76> / cell_PIM
XI21767 bl<56> cbl<28> in1<99> in2<99> sl<56> vdd vss wl<99> / cell_PIM
XI21766 bl<56> cbl<28> in1<100> in2<100> sl<56> vdd vss wl<100> / cell_PIM
XI21765 bl<56> cbl<28> in1<102> in2<102> sl<56> vdd vss wl<102> / cell_PIM
XI21764 bl<56> cbl<28> in1<103> in2<103> sl<56> vdd vss wl<103> / cell_PIM
XI21118 bl<48> cbl<24> in1<118> in2<118> sl<48> vdd vss wl<118> / cell_PIM
XI21117 bl<48> cbl<24> in1<122> in2<122> sl<48> vdd vss wl<122> / cell_PIM
XI21116 bl<48> cbl<24> in1<121> in2<121> sl<48> vdd vss wl<121> / cell_PIM
XI21115 bl<48> cbl<24> in1<120> in2<120> sl<48> vdd vss wl<120> / cell_PIM
XI22414 bl<32> cbl<16> in1<75> in2<75> sl<32> vdd vss wl<75> / cell_PIM
XI21109 bl<46> cbl<23> in1<118> in2<118> sl<46> vdd vss wl<118> / cell_PIM
XI21763 bl<56> cbl<28> in1<101> in2<101> sl<56> vdd vss wl<101> / cell_PIM
XI22412 bl<32> cbl<16> in1<78> in2<78> sl<32> vdd vss wl<78> / cell_PIM
XI22411 bl<32> cbl<16> in1<77> in2<77> sl<32> vdd vss wl<77> / cell_PIM
XI21108 bl<46> cbl<23> in1<119> in2<119> sl<46> vdd vss wl<119> / cell_PIM
XI21107 bl<46> cbl<23> in1<121> in2<121> sl<46> vdd vss wl<121> / cell_PIM
XI21106 bl<46> cbl<23> in1<122> in2<122> sl<46> vdd vss wl<122> / cell_PIM
XI21105 bl<46> cbl<23> in1<120> in2<120> sl<46> vdd vss wl<120> / cell_PIM
XI21757 bl<54> cbl<27> in1<99> in2<99> sl<54> vdd vss wl<99> / cell_PIM
XI21756 bl<54> cbl<27> in1<100> in2<100> sl<54> vdd vss wl<100> / cell_PIM
XI21755 bl<54> cbl<27> in1<102> in2<102> sl<54> vdd vss wl<102> / cell_PIM
XI21754 bl<54> cbl<27> in1<103> in2<103> sl<54> vdd vss wl<103> / cell_PIM
XI22406 bl<62> cbl<31> in1<80> in2<80> sl<62> vdd vss wl<80> / cell_PIM
XI22405 bl<62> cbl<31> in1<81> in2<81> sl<62> vdd vss wl<81> / cell_PIM
XI22404 bl<62> cbl<31> in1<83> in2<83> sl<62> vdd vss wl<83> / cell_PIM
XI19442 bl<30> cbl<15> in1<93> in2<93> sl<30> vdd vss wl<93> / cell_PIM
XI19441 bl<30> cbl<15> in1<92> in2<92> sl<30> vdd vss wl<92> / cell_PIM
XI19443 bl<30> cbl<15> in1<91> in2<91> sl<30> vdd vss wl<91> / cell_PIM
XI20611 bl<20> cbl<10> in1<14> in2<14> sl<20> vdd vss wl<14> / cell_PIM
XI20610 bl<20> cbl<10> in1<13> in2<13> sl<20> vdd vss wl<13> / cell_PIM
XI20609 bl<20> cbl<10> in1<17> in2<17> sl<20> vdd vss wl<17> / cell_PIM
XI20608 bl<20> cbl<10> in1<16> in2<16> sl<20> vdd vss wl<16> / cell_PIM
XI20607 bl<20> cbl<10> in1<15> in2<15> sl<20> vdd vss wl<15> / cell_PIM
XI20023 bl<24> cbl<12> in1<51> in2<51> sl<24> vdd vss wl<51> / cell_PIM
XI20022 bl<24> cbl<12> in1<52> in2<52> sl<24> vdd vss wl<52> / cell_PIM
XI20021 bl<24> cbl<12> in1<54> in2<54> sl<24> vdd vss wl<54> / cell_PIM
XI19435 bl<28> cbl<14> in1<91> in2<91> sl<28> vdd vss wl<91> / cell_PIM
XI19434 bl<28> cbl<14> in1<90> in2<90> sl<28> vdd vss wl<90> / cell_PIM
XI19432 bl<28> cbl<14> in1<93> in2<93> sl<28> vdd vss wl<93> / cell_PIM
XI19431 bl<28> cbl<14> in1<92> in2<92> sl<28> vdd vss wl<92> / cell_PIM
XI19433 bl<28> cbl<14> in1<89> in2<89> sl<28> vdd vss wl<89> / cell_PIM
XI20020 bl<24> cbl<12> in1<55> in2<55> sl<24> vdd vss wl<55> / cell_PIM
XI20019 bl<24> cbl<12> in1<53> in2<53> sl<24> vdd vss wl<53> / cell_PIM
XI20601 bl<18> cbl<9> in1<13> in2<13> sl<18> vdd vss wl<13> / cell_PIM
XI20600 bl<18> cbl<9> in1<14> in2<14> sl<18> vdd vss wl<14> / cell_PIM
XI20599 bl<18> cbl<9> in1<16> in2<16> sl<18> vdd vss wl<16> / cell_PIM
XI19425 bl<26> cbl<13> in1<89> in2<89> sl<26> vdd vss wl<89> / cell_PIM
XI19424 bl<26> cbl<13> in1<90> in2<90> sl<26> vdd vss wl<90> / cell_PIM
XI20013 bl<22> cbl<11> in1<51> in2<51> sl<22> vdd vss wl<51> / cell_PIM
XI20598 bl<18> cbl<9> in1<17> in2<17> sl<18> vdd vss wl<17> / cell_PIM
XI20597 bl<18> cbl<9> in1<15> in2<15> sl<18> vdd vss wl<15> / cell_PIM
XI19422 bl<26> cbl<13> in1<93> in2<93> sl<26> vdd vss wl<93> / cell_PIM
XI19421 bl<26> cbl<13> in1<92> in2<92> sl<26> vdd vss wl<92> / cell_PIM
XI19423 bl<26> cbl<13> in1<91> in2<91> sl<26> vdd vss wl<91> / cell_PIM
XI20012 bl<22> cbl<11> in1<52> in2<52> sl<22> vdd vss wl<52> / cell_PIM
XI20011 bl<22> cbl<11> in1<54> in2<54> sl<22> vdd vss wl<54> / cell_PIM
XI20010 bl<22> cbl<11> in1<55> in2<55> sl<22> vdd vss wl<55> / cell_PIM
XI20009 bl<22> cbl<11> in1<53> in2<53> sl<22> vdd vss wl<53> / cell_PIM
XI20591 bl<16> cbl<8> in1<14> in2<14> sl<16> vdd vss wl<14> / cell_PIM
XI20590 bl<16> cbl<8> in1<13> in2<13> sl<16> vdd vss wl<13> / cell_PIM
XI20589 bl<16> cbl<8> in1<17> in2<17> sl<16> vdd vss wl<17> / cell_PIM
XI20588 bl<16> cbl<8> in1<16> in2<16> sl<16> vdd vss wl<16> / cell_PIM
XI20587 bl<16> cbl<8> in1<15> in2<15> sl<16> vdd vss wl<15> / cell_PIM
XI19415 bl<24> cbl<12> in1<89> in2<89> sl<24> vdd vss wl<89> / cell_PIM
XI19414 bl<24> cbl<12> in1<90> in2<90> sl<24> vdd vss wl<90> / cell_PIM
XI19412 bl<24> cbl<12> in1<93> in2<93> sl<24> vdd vss wl<93> / cell_PIM
XI19411 bl<24> cbl<12> in1<92> in2<92> sl<24> vdd vss wl<92> / cell_PIM
XI19413 bl<24> cbl<12> in1<91> in2<91> sl<24> vdd vss wl<91> / cell_PIM
XI20003 bl<20> cbl<10> in1<52> in2<52> sl<20> vdd vss wl<52> / cell_PIM
XI20002 bl<20> cbl<10> in1<51> in2<51> sl<20> vdd vss wl<51> / cell_PIM
XI20001 bl<20> cbl<10> in1<55> in2<55> sl<20> vdd vss wl<55> / cell_PIM
XI20582 bl<30> cbl<15> in1<18> in2<18> sl<30> vdd vss wl<18> / cell_PIM
XI20581 bl<30> cbl<15> in1<19> in2<19> sl<30> vdd vss wl<19> / cell_PIM
XI20580 bl<30> cbl<15> in1<21> in2<21> sl<30> vdd vss wl<21> / cell_PIM
XI20579 bl<30> cbl<15> in1<20> in2<20> sl<30> vdd vss wl<20> / cell_PIM
XI19405 bl<22> cbl<11> in1<89> in2<89> sl<22> vdd vss wl<89> / cell_PIM
XI19404 bl<22> cbl<11> in1<90> in2<90> sl<22> vdd vss wl<90> / cell_PIM
XI20000 bl<20> cbl<10> in1<54> in2<54> sl<20> vdd vss wl<54> / cell_PIM
XI19999 bl<20> cbl<10> in1<53> in2<53> sl<20> vdd vss wl<53> / cell_PIM
XI20574 bl<28> cbl<14> in1<19> in2<19> sl<28> vdd vss wl<19> / cell_PIM
XI19402 bl<22> cbl<11> in1<93> in2<93> sl<22> vdd vss wl<93> / cell_PIM
XI19401 bl<22> cbl<11> in1<92> in2<92> sl<22> vdd vss wl<92> / cell_PIM
XI19403 bl<22> cbl<11> in1<91> in2<91> sl<22> vdd vss wl<91> / cell_PIM
XI19993 bl<18> cbl<9> in1<51> in2<51> sl<18> vdd vss wl<51> / cell_PIM
XI20573 bl<28> cbl<14> in1<18> in2<18> sl<28> vdd vss wl<18> / cell_PIM
XI20572 bl<28> cbl<14> in1<21> in2<21> sl<28> vdd vss wl<21> / cell_PIM
XI20571 bl<28> cbl<14> in1<20> in2<20> sl<28> vdd vss wl<20> / cell_PIM
XI20566 bl<26> cbl<13> in1<18> in2<18> sl<26> vdd vss wl<18> / cell_PIM
XI20565 bl<26> cbl<13> in1<19> in2<19> sl<26> vdd vss wl<19> / cell_PIM
XI20564 bl<26> cbl<13> in1<21> in2<21> sl<26> vdd vss wl<21> / cell_PIM
XI19992 bl<18> cbl<9> in1<52> in2<52> sl<18> vdd vss wl<52> / cell_PIM
XI19991 bl<18> cbl<9> in1<54> in2<54> sl<18> vdd vss wl<54> / cell_PIM
XI19990 bl<18> cbl<9> in1<55> in2<55> sl<18> vdd vss wl<55> / cell_PIM
XI19989 bl<18> cbl<9> in1<53> in2<53> sl<18> vdd vss wl<53> / cell_PIM
XI19395 bl<20> cbl<10> in1<91> in2<91> sl<20> vdd vss wl<91> / cell_PIM
XI19394 bl<20> cbl<10> in1<90> in2<90> sl<20> vdd vss wl<90> / cell_PIM
XI19392 bl<20> cbl<10> in1<93> in2<93> sl<20> vdd vss wl<93> / cell_PIM
XI19391 bl<20> cbl<10> in1<92> in2<92> sl<20> vdd vss wl<92> / cell_PIM
XI19393 bl<20> cbl<10> in1<89> in2<89> sl<20> vdd vss wl<89> / cell_PIM
XI20563 bl<26> cbl<13> in1<20> in2<20> sl<26> vdd vss wl<20> / cell_PIM
XI19385 bl<18> cbl<9> in1<89> in2<89> sl<18> vdd vss wl<89> / cell_PIM
XI19384 bl<18> cbl<9> in1<90> in2<90> sl<18> vdd vss wl<90> / cell_PIM
XI19983 bl<16> cbl<8> in1<52> in2<52> sl<16> vdd vss wl<52> / cell_PIM
XI19982 bl<16> cbl<8> in1<51> in2<51> sl<16> vdd vss wl<51> / cell_PIM
XI19981 bl<16> cbl<8> in1<55> in2<55> sl<16> vdd vss wl<55> / cell_PIM
XI20558 bl<24> cbl<12> in1<18> in2<18> sl<24> vdd vss wl<18> / cell_PIM
XI20557 bl<24> cbl<12> in1<19> in2<19> sl<24> vdd vss wl<19> / cell_PIM
XI20556 bl<24> cbl<12> in1<21> in2<21> sl<24> vdd vss wl<21> / cell_PIM
XI20555 bl<24> cbl<12> in1<20> in2<20> sl<24> vdd vss wl<20> / cell_PIM
XI19382 bl<18> cbl<9> in1<93> in2<93> sl<18> vdd vss wl<93> / cell_PIM
XI19381 bl<18> cbl<9> in1<92> in2<92> sl<18> vdd vss wl<92> / cell_PIM
XI19383 bl<18> cbl<9> in1<91> in2<91> sl<18> vdd vss wl<91> / cell_PIM
XI19980 bl<16> cbl<8> in1<54> in2<54> sl<16> vdd vss wl<54> / cell_PIM
XI19979 bl<16> cbl<8> in1<53> in2<53> sl<16> vdd vss wl<53> / cell_PIM
XI20550 bl<22> cbl<11> in1<18> in2<18> sl<22> vdd vss wl<18> / cell_PIM
XI20549 bl<22> cbl<11> in1<19> in2<19> sl<22> vdd vss wl<19> / cell_PIM
XI20548 bl<22> cbl<11> in1<21> in2<21> sl<22> vdd vss wl<21> / cell_PIM
XI20547 bl<22> cbl<11> in1<20> in2<20> sl<22> vdd vss wl<20> / cell_PIM
XI19973 bl<30> cbl<15> in1<56> in2<56> sl<30> vdd vss wl<56> / cell_PIM
XI19375 bl<16> cbl<8> in1<91> in2<91> sl<16> vdd vss wl<91> / cell_PIM
XI19374 bl<16> cbl<8> in1<90> in2<90> sl<16> vdd vss wl<90> / cell_PIM
XI19372 bl<16> cbl<8> in1<93> in2<93> sl<16> vdd vss wl<93> / cell_PIM
XI19371 bl<16> cbl<8> in1<92> in2<92> sl<16> vdd vss wl<92> / cell_PIM
XI19373 bl<16> cbl<8> in1<89> in2<89> sl<16> vdd vss wl<89> / cell_PIM
XI19972 bl<30> cbl<15> in1<57> in2<57> sl<30> vdd vss wl<57> / cell_PIM
XI19971 bl<30> cbl<15> in1<59> in2<59> sl<30> vdd vss wl<59> / cell_PIM
XI19970 bl<30> cbl<15> in1<60> in2<60> sl<30> vdd vss wl<60> / cell_PIM
XI19969 bl<30> cbl<15> in1<58> in2<58> sl<30> vdd vss wl<58> / cell_PIM
XI20542 bl<20> cbl<10> in1<19> in2<19> sl<20> vdd vss wl<19> / cell_PIM
XI20541 bl<20> cbl<10> in1<18> in2<18> sl<20> vdd vss wl<18> / cell_PIM
XI20540 bl<20> cbl<10> in1<21> in2<21> sl<20> vdd vss wl<21> / cell_PIM
XI20539 bl<20> cbl<10> in1<20> in2<20> sl<20> vdd vss wl<20> / cell_PIM
XI19365 bl<30> cbl<15> in1<94> in2<94> sl<30> vdd vss wl<94> / cell_PIM
XI19364 bl<30> cbl<15> in1<95> in2<95> sl<30> vdd vss wl<95> / cell_PIM
XI20534 bl<18> cbl<9> in1<18> in2<18> sl<18> vdd vss wl<18> / cell_PIM
XI19362 bl<30> cbl<15> in1<98> in2<98> sl<30> vdd vss wl<98> / cell_PIM
XI19361 bl<30> cbl<15> in1<96> in2<96> sl<30> vdd vss wl<96> / cell_PIM
XI19363 bl<30> cbl<15> in1<97> in2<97> sl<30> vdd vss wl<97> / cell_PIM
XI19963 bl<28> cbl<14> in1<57> in2<57> sl<28> vdd vss wl<57> / cell_PIM
XI19962 bl<28> cbl<14> in1<56> in2<56> sl<28> vdd vss wl<56> / cell_PIM
XI19961 bl<28> cbl<14> in1<60> in2<60> sl<28> vdd vss wl<60> / cell_PIM
XI20533 bl<18> cbl<9> in1<19> in2<19> sl<18> vdd vss wl<19> / cell_PIM
XI20532 bl<18> cbl<9> in1<21> in2<21> sl<18> vdd vss wl<21> / cell_PIM
XI20531 bl<18> cbl<9> in1<20> in2<20> sl<18> vdd vss wl<20> / cell_PIM
XI20526 bl<16> cbl<8> in1<19> in2<19> sl<16> vdd vss wl<19> / cell_PIM
XI20525 bl<16> cbl<8> in1<18> in2<18> sl<16> vdd vss wl<18> / cell_PIM
XI20524 bl<16> cbl<8> in1<21> in2<21> sl<16> vdd vss wl<21> / cell_PIM
XI19960 bl<28> cbl<14> in1<59> in2<59> sl<28> vdd vss wl<59> / cell_PIM
XI19959 bl<28> cbl<14> in1<58> in2<58> sl<28> vdd vss wl<58> / cell_PIM
XI19355 bl<28> cbl<14> in1<95> in2<95> sl<28> vdd vss wl<95> / cell_PIM
XI19354 bl<28> cbl<14> in1<94> in2<94> sl<28> vdd vss wl<94> / cell_PIM
XI19352 bl<28> cbl<14> in1<97> in2<97> sl<28> vdd vss wl<97> / cell_PIM
XI19351 bl<28> cbl<14> in1<96> in2<96> sl<28> vdd vss wl<96> / cell_PIM
XI19353 bl<28> cbl<14> in1<98> in2<98> sl<28> vdd vss wl<98> / cell_PIM
XI19953 bl<26> cbl<13> in1<56> in2<56> sl<26> vdd vss wl<56> / cell_PIM
XI20523 bl<16> cbl<8> in1<20> in2<20> sl<16> vdd vss wl<20> / cell_PIM
XI19345 bl<26> cbl<13> in1<94> in2<94> sl<26> vdd vss wl<94> / cell_PIM
XI19344 bl<26> cbl<13> in1<95> in2<95> sl<26> vdd vss wl<95> / cell_PIM
XI19952 bl<26> cbl<13> in1<57> in2<57> sl<26> vdd vss wl<57> / cell_PIM
XI19951 bl<26> cbl<13> in1<59> in2<59> sl<26> vdd vss wl<59> / cell_PIM
XI19950 bl<26> cbl<13> in1<60> in2<60> sl<26> vdd vss wl<60> / cell_PIM
XI19949 bl<26> cbl<13> in1<58> in2<58> sl<26> vdd vss wl<58> / cell_PIM
XI20517 bl<30> cbl<15> in1<22> in2<22> sl<30> vdd vss wl<22> / cell_PIM
XI20516 bl<30> cbl<15> in1<23> in2<23> sl<30> vdd vss wl<23> / cell_PIM
XI20515 bl<30> cbl<15> in1<24> in2<24> sl<30> vdd vss wl<24> / cell_PIM
XI20514 bl<30> cbl<15> in1<26> in2<26> sl<30> vdd vss wl<26> / cell_PIM
XI19342 bl<26> cbl<13> in1<98> in2<98> sl<26> vdd vss wl<98> / cell_PIM
XI19341 bl<26> cbl<13> in1<96> in2<96> sl<26> vdd vss wl<96> / cell_PIM
XI19343 bl<26> cbl<13> in1<97> in2<97> sl<26> vdd vss wl<97> / cell_PIM
XI20513 bl<30> cbl<15> in1<25> in2<25> sl<30> vdd vss wl<25> / cell_PIM
XI20507 bl<28> cbl<14> in1<24> in2<24> sl<28> vdd vss wl<24> / cell_PIM
XI20506 bl<28> cbl<14> in1<23> in2<23> sl<28> vdd vss wl<23> / cell_PIM
XI20505 bl<28> cbl<14> in1<22> in2<22> sl<28> vdd vss wl<22> / cell_PIM
XI20504 bl<28> cbl<14> in1<26> in2<26> sl<28> vdd vss wl<26> / cell_PIM
XI19943 bl<24> cbl<12> in1<56> in2<56> sl<24> vdd vss wl<56> / cell_PIM
XI19942 bl<24> cbl<12> in1<57> in2<57> sl<24> vdd vss wl<57> / cell_PIM
XI19941 bl<24> cbl<12> in1<59> in2<59> sl<24> vdd vss wl<59> / cell_PIM
XI19335 bl<24> cbl<12> in1<94> in2<94> sl<24> vdd vss wl<94> / cell_PIM
XI19334 bl<24> cbl<12> in1<95> in2<95> sl<24> vdd vss wl<95> / cell_PIM
XI19332 bl<24> cbl<12> in1<98> in2<98> sl<24> vdd vss wl<98> / cell_PIM
XI19331 bl<24> cbl<12> in1<96> in2<96> sl<24> vdd vss wl<96> / cell_PIM
XI19333 bl<24> cbl<12> in1<97> in2<97> sl<24> vdd vss wl<97> / cell_PIM
XI19940 bl<24> cbl<12> in1<60> in2<60> sl<24> vdd vss wl<60> / cell_PIM
XI19939 bl<24> cbl<12> in1<58> in2<58> sl<24> vdd vss wl<58> / cell_PIM
XI20503 bl<28> cbl<14> in1<25> in2<25> sl<28> vdd vss wl<25> / cell_PIM
XI19325 bl<22> cbl<11> in1<94> in2<94> sl<22> vdd vss wl<94> / cell_PIM
XI19324 bl<22> cbl<11> in1<95> in2<95> sl<22> vdd vss wl<95> / cell_PIM
XI19933 bl<22> cbl<11> in1<56> in2<56> sl<22> vdd vss wl<56> / cell_PIM
XI20497 bl<26> cbl<13> in1<22> in2<22> sl<26> vdd vss wl<22> / cell_PIM
XI20496 bl<26> cbl<13> in1<23> in2<23> sl<26> vdd vss wl<23> / cell_PIM
XI20495 bl<26> cbl<13> in1<24> in2<24> sl<26> vdd vss wl<24> / cell_PIM
XI20494 bl<26> cbl<13> in1<26> in2<26> sl<26> vdd vss wl<26> / cell_PIM
XI19322 bl<22> cbl<11> in1<98> in2<98> sl<22> vdd vss wl<98> / cell_PIM
XI19321 bl<22> cbl<11> in1<96> in2<96> sl<22> vdd vss wl<96> / cell_PIM
XI19323 bl<22> cbl<11> in1<97> in2<97> sl<22> vdd vss wl<97> / cell_PIM
XI19932 bl<22> cbl<11> in1<57> in2<57> sl<22> vdd vss wl<57> / cell_PIM
XI19931 bl<22> cbl<11> in1<59> in2<59> sl<22> vdd vss wl<59> / cell_PIM
XI19930 bl<22> cbl<11> in1<60> in2<60> sl<22> vdd vss wl<60> / cell_PIM
XI19929 bl<22> cbl<11> in1<58> in2<58> sl<22> vdd vss wl<58> / cell_PIM
XI20493 bl<26> cbl<13> in1<25> in2<25> sl<26> vdd vss wl<25> / cell_PIM
XI20487 bl<24> cbl<12> in1<22> in2<22> sl<24> vdd vss wl<22> / cell_PIM
XI20486 bl<24> cbl<12> in1<23> in2<23> sl<24> vdd vss wl<23> / cell_PIM
XI20485 bl<24> cbl<12> in1<24> in2<24> sl<24> vdd vss wl<24> / cell_PIM
XI20484 bl<24> cbl<12> in1<26> in2<26> sl<24> vdd vss wl<26> / cell_PIM
XI19315 bl<20> cbl<10> in1<95> in2<95> sl<20> vdd vss wl<95> / cell_PIM
XI19314 bl<20> cbl<10> in1<94> in2<94> sl<20> vdd vss wl<94> / cell_PIM
XI19312 bl<20> cbl<10> in1<97> in2<97> sl<20> vdd vss wl<97> / cell_PIM
XI19311 bl<20> cbl<10> in1<96> in2<96> sl<20> vdd vss wl<96> / cell_PIM
XI19313 bl<20> cbl<10> in1<98> in2<98> sl<20> vdd vss wl<98> / cell_PIM
XI19923 bl<20> cbl<10> in1<57> in2<57> sl<20> vdd vss wl<57> / cell_PIM
XI19922 bl<20> cbl<10> in1<56> in2<56> sl<20> vdd vss wl<56> / cell_PIM
XI19921 bl<20> cbl<10> in1<60> in2<60> sl<20> vdd vss wl<60> / cell_PIM
XI20483 bl<24> cbl<12> in1<25> in2<25> sl<24> vdd vss wl<25> / cell_PIM
XI19305 bl<18> cbl<9> in1<94> in2<94> sl<18> vdd vss wl<94> / cell_PIM
XI19304 bl<18> cbl<9> in1<95> in2<95> sl<18> vdd vss wl<95> / cell_PIM
XI19920 bl<20> cbl<10> in1<59> in2<59> sl<20> vdd vss wl<59> / cell_PIM
XI19919 bl<20> cbl<10> in1<58> in2<58> sl<20> vdd vss wl<58> / cell_PIM
XI20477 bl<22> cbl<11> in1<22> in2<22> sl<22> vdd vss wl<22> / cell_PIM
XI20476 bl<22> cbl<11> in1<23> in2<23> sl<22> vdd vss wl<23> / cell_PIM
XI20475 bl<22> cbl<11> in1<24> in2<24> sl<22> vdd vss wl<24> / cell_PIM
XI20474 bl<22> cbl<11> in1<26> in2<26> sl<22> vdd vss wl<26> / cell_PIM
XI19302 bl<18> cbl<9> in1<98> in2<98> sl<18> vdd vss wl<98> / cell_PIM
XI19301 bl<18> cbl<9> in1<96> in2<96> sl<18> vdd vss wl<96> / cell_PIM
XI19303 bl<18> cbl<9> in1<97> in2<97> sl<18> vdd vss wl<97> / cell_PIM
XI19913 bl<18> cbl<9> in1<56> in2<56> sl<18> vdd vss wl<56> / cell_PIM
XI20473 bl<22> cbl<11> in1<25> in2<25> sl<22> vdd vss wl<25> / cell_PIM
XI20467 bl<20> cbl<10> in1<24> in2<24> sl<20> vdd vss wl<24> / cell_PIM
XI20466 bl<20> cbl<10> in1<23> in2<23> sl<20> vdd vss wl<23> / cell_PIM
XI20465 bl<20> cbl<10> in1<22> in2<22> sl<20> vdd vss wl<22> / cell_PIM
XI20464 bl<20> cbl<10> in1<26> in2<26> sl<20> vdd vss wl<26> / cell_PIM
XI19912 bl<18> cbl<9> in1<57> in2<57> sl<18> vdd vss wl<57> / cell_PIM
XI19911 bl<18> cbl<9> in1<59> in2<59> sl<18> vdd vss wl<59> / cell_PIM
XI19910 bl<18> cbl<9> in1<60> in2<60> sl<18> vdd vss wl<60> / cell_PIM
XI19909 bl<18> cbl<9> in1<58> in2<58> sl<18> vdd vss wl<58> / cell_PIM
XI19295 bl<16> cbl<8> in1<95> in2<95> sl<16> vdd vss wl<95> / cell_PIM
XI19294 bl<16> cbl<8> in1<94> in2<94> sl<16> vdd vss wl<94> / cell_PIM
XI19292 bl<16> cbl<8> in1<97> in2<97> sl<16> vdd vss wl<97> / cell_PIM
XI19291 bl<16> cbl<8> in1<96> in2<96> sl<16> vdd vss wl<96> / cell_PIM
XI19293 bl<16> cbl<8> in1<98> in2<98> sl<16> vdd vss wl<98> / cell_PIM
XI20463 bl<20> cbl<10> in1<25> in2<25> sl<20> vdd vss wl<25> / cell_PIM
XI19285 bl<30> cbl<15> in1<99> in2<99> sl<30> vdd vss wl<99> / cell_PIM
XI19284 bl<30> cbl<15> in1<100> in2<100> sl<30> vdd vss wl<100> / cell_PIM
XI19903 bl<16> cbl<8> in1<57> in2<57> sl<16> vdd vss wl<57> / cell_PIM
XI19902 bl<16> cbl<8> in1<56> in2<56> sl<16> vdd vss wl<56> / cell_PIM
XI19901 bl<16> cbl<8> in1<60> in2<60> sl<16> vdd vss wl<60> / cell_PIM
XI20457 bl<18> cbl<9> in1<22> in2<22> sl<18> vdd vss wl<22> / cell_PIM
XI20456 bl<18> cbl<9> in1<23> in2<23> sl<18> vdd vss wl<23> / cell_PIM
XI20455 bl<18> cbl<9> in1<24> in2<24> sl<18> vdd vss wl<24> / cell_PIM
XI20454 bl<18> cbl<9> in1<26> in2<26> sl<18> vdd vss wl<26> / cell_PIM
XI17489 bl<6> cbl<3> in1<78> in2<78> sl<6> vdd vss wl<78> / cell_PIM
XI18143 bl<10> cbl<5> in1<85> in2<85> sl<10> vdd vss wl<85> / cell_PIM
XI18142 bl<10> cbl<5> in1<86> in2<86> sl<10> vdd vss wl<86> / cell_PIM
XI18141 bl<10> cbl<5> in1<82> in2<82> sl<10> vdd vss wl<82> / cell_PIM
XI18790 bl<8> cbl<4> in1<4> in2<4> sl<8> vdd vss wl<4> / cell_PIM
XI18789 bl<8> cbl<4> in1<3> in2<3> sl<8> vdd vss wl<3> / cell_PIM
XI18788 bl<8> cbl<4> in1<2> in2<2> sl<8> vdd vss wl<2> / cell_PIM
XI18787 bl<8> cbl<4> in1<1> in2<1> sl<8> vdd vss wl<1> / cell_PIM
XI18135 bl<8> cbl<4> in1<86> in2<86> sl<8> vdd vss wl<86> / cell_PIM
XI18134 bl<8> cbl<4> in1<85> in2<85> sl<8> vdd vss wl<85> / cell_PIM
XI17488 bl<6> cbl<3> in1<79> in2<79> sl<6> vdd vss wl<79> / cell_PIM
XI17487 bl<6> cbl<3> in1<80> in2<80> sl<6> vdd vss wl<80> / cell_PIM
XI17486 bl<6> cbl<3> in1<81> in2<81> sl<6> vdd vss wl<81> / cell_PIM
XI17485 bl<6> cbl<3> in1<77> in2<77> sl<6> vdd vss wl<77> / cell_PIM
XI17479 bl<4> cbl<2> in1<81> in2<81> sl<4> vdd vss wl<81> / cell_PIM
XI18133 bl<8> cbl<4> in1<84> in2<84> sl<8> vdd vss wl<84> / cell_PIM
XI18132 bl<8> cbl<4> in1<83> in2<83> sl<8> vdd vss wl<83> / cell_PIM
XI18131 bl<8> cbl<4> in1<82> in2<82> sl<8> vdd vss wl<82> / cell_PIM
XI18781 bl<14> cbl<7> in1<6> in2<6> sl<14> vdd vss wl<6> / cell_PIM
XI18780 bl<14> cbl<7> in1<7> in2<7> sl<14> vdd vss wl<7> / cell_PIM
XI18779 bl<14> cbl<7> in1<8> in2<8> sl<14> vdd vss wl<8> / cell_PIM
XI17478 bl<4> cbl<2> in1<80> in2<80> sl<4> vdd vss wl<80> / cell_PIM
XI17477 bl<4> cbl<2> in1<79> in2<79> sl<4> vdd vss wl<79> / cell_PIM
XI17476 bl<4> cbl<2> in1<78> in2<78> sl<4> vdd vss wl<78> / cell_PIM
XI17475 bl<4> cbl<2> in1<77> in2<77> sl<4> vdd vss wl<77> / cell_PIM
XI18125 bl<14> cbl<7> in1<88> in2<88> sl<14> vdd vss wl<88> / cell_PIM
XI18124 bl<14> cbl<7> in1<89> in2<89> sl<14> vdd vss wl<89> / cell_PIM
XI18778 bl<14> cbl<7> in1<9> in2<9> sl<14> vdd vss wl<9> / cell_PIM
XI18777 bl<14> cbl<7> in1<5> in2<5> sl<14> vdd vss wl<5> / cell_PIM
XI17469 bl<6> cbl<3> in1<83> in2<83> sl<6> vdd vss wl<83> / cell_PIM
XI18123 bl<14> cbl<7> in1<90> in2<90> sl<14> vdd vss wl<90> / cell_PIM
XI18122 bl<14> cbl<7> in1<91> in2<91> sl<14> vdd vss wl<91> / cell_PIM
XI18121 bl<14> cbl<7> in1<87> in2<87> sl<14> vdd vss wl<87> / cell_PIM
XI18771 bl<12> cbl<6> in1<9> in2<9> sl<12> vdd vss wl<9> / cell_PIM
XI18770 bl<12> cbl<6> in1<8> in2<8> sl<12> vdd vss wl<8> / cell_PIM
XI18769 bl<12> cbl<6> in1<7> in2<7> sl<12> vdd vss wl<7> / cell_PIM
XI18768 bl<12> cbl<6> in1<6> in2<6> sl<12> vdd vss wl<6> / cell_PIM
XI18767 bl<12> cbl<6> in1<5> in2<5> sl<12> vdd vss wl<5> / cell_PIM
XI18115 bl<12> cbl<6> in1<91> in2<91> sl<12> vdd vss wl<91> / cell_PIM
XI18114 bl<12> cbl<6> in1<90> in2<90> sl<12> vdd vss wl<90> / cell_PIM
XI17468 bl<6> cbl<3> in1<84> in2<84> sl<6> vdd vss wl<84> / cell_PIM
XI17467 bl<6> cbl<3> in1<85> in2<85> sl<6> vdd vss wl<85> / cell_PIM
XI17466 bl<6> cbl<3> in1<86> in2<86> sl<6> vdd vss wl<86> / cell_PIM
XI17465 bl<6> cbl<3> in1<82> in2<82> sl<6> vdd vss wl<82> / cell_PIM
XI17459 bl<4> cbl<2> in1<86> in2<86> sl<4> vdd vss wl<86> / cell_PIM
XI18113 bl<12> cbl<6> in1<89> in2<89> sl<12> vdd vss wl<89> / cell_PIM
XI18112 bl<12> cbl<6> in1<88> in2<88> sl<12> vdd vss wl<88> / cell_PIM
XI18111 bl<12> cbl<6> in1<87> in2<87> sl<12> vdd vss wl<87> / cell_PIM
XI18761 bl<10> cbl<5> in1<6> in2<6> sl<10> vdd vss wl<6> / cell_PIM
XI18760 bl<10> cbl<5> in1<7> in2<7> sl<10> vdd vss wl<7> / cell_PIM
XI18759 bl<10> cbl<5> in1<8> in2<8> sl<10> vdd vss wl<8> / cell_PIM
XI17458 bl<4> cbl<2> in1<85> in2<85> sl<4> vdd vss wl<85> / cell_PIM
XI17457 bl<4> cbl<2> in1<84> in2<84> sl<4> vdd vss wl<84> / cell_PIM
XI17456 bl<4> cbl<2> in1<83> in2<83> sl<4> vdd vss wl<83> / cell_PIM
XI17455 bl<4> cbl<2> in1<82> in2<82> sl<4> vdd vss wl<82> / cell_PIM
XI18105 bl<10> cbl<5> in1<88> in2<88> sl<10> vdd vss wl<88> / cell_PIM
XI18104 bl<10> cbl<5> in1<89> in2<89> sl<10> vdd vss wl<89> / cell_PIM
XI18758 bl<10> cbl<5> in1<9> in2<9> sl<10> vdd vss wl<9> / cell_PIM
XI18757 bl<10> cbl<5> in1<5> in2<5> sl<10> vdd vss wl<5> / cell_PIM
XI17449 bl<6> cbl<3> in1<88> in2<88> sl<6> vdd vss wl<88> / cell_PIM
XI18103 bl<10> cbl<5> in1<90> in2<90> sl<10> vdd vss wl<90> / cell_PIM
XI18102 bl<10> cbl<5> in1<91> in2<91> sl<10> vdd vss wl<91> / cell_PIM
XI18101 bl<10> cbl<5> in1<87> in2<87> sl<10> vdd vss wl<87> / cell_PIM
XI18751 bl<8> cbl<4> in1<9> in2<9> sl<8> vdd vss wl<9> / cell_PIM
XI18750 bl<8> cbl<4> in1<8> in2<8> sl<8> vdd vss wl<8> / cell_PIM
XI18749 bl<8> cbl<4> in1<7> in2<7> sl<8> vdd vss wl<7> / cell_PIM
XI18748 bl<8> cbl<4> in1<6> in2<6> sl<8> vdd vss wl<6> / cell_PIM
XI18747 bl<8> cbl<4> in1<5> in2<5> sl<8> vdd vss wl<5> / cell_PIM
XI18095 bl<8> cbl<4> in1<91> in2<91> sl<8> vdd vss wl<91> / cell_PIM
XI18094 bl<8> cbl<4> in1<90> in2<90> sl<8> vdd vss wl<90> / cell_PIM
XI17448 bl<6> cbl<3> in1<89> in2<89> sl<6> vdd vss wl<89> / cell_PIM
XI17447 bl<6> cbl<3> in1<90> in2<90> sl<6> vdd vss wl<90> / cell_PIM
XI17446 bl<6> cbl<3> in1<91> in2<91> sl<6> vdd vss wl<91> / cell_PIM
XI17445 bl<6> cbl<3> in1<87> in2<87> sl<6> vdd vss wl<87> / cell_PIM
XI17439 bl<4> cbl<2> in1<91> in2<91> sl<4> vdd vss wl<91> / cell_PIM
XI18093 bl<8> cbl<4> in1<89> in2<89> sl<8> vdd vss wl<89> / cell_PIM
XI18092 bl<8> cbl<4> in1<88> in2<88> sl<8> vdd vss wl<88> / cell_PIM
XI18091 bl<8> cbl<4> in1<87> in2<87> sl<8> vdd vss wl<87> / cell_PIM
XI18741 bl<14> cbl<7> in1<11> in2<11> sl<14> vdd vss wl<11> / cell_PIM
XI18740 bl<14> cbl<7> in1<12> in2<12> sl<14> vdd vss wl<12> / cell_PIM
XI18739 bl<14> cbl<7> in1<13> in2<13> sl<14> vdd vss wl<13> / cell_PIM
XI17438 bl<4> cbl<2> in1<90> in2<90> sl<4> vdd vss wl<90> / cell_PIM
XI17437 bl<4> cbl<2> in1<89> in2<89> sl<4> vdd vss wl<89> / cell_PIM
XI17436 bl<4> cbl<2> in1<88> in2<88> sl<4> vdd vss wl<88> / cell_PIM
XI17435 bl<4> cbl<2> in1<87> in2<87> sl<4> vdd vss wl<87> / cell_PIM
XI18086 bl<14> cbl<7> in1<93> in2<93> sl<14> vdd vss wl<93> / cell_PIM
XI18085 bl<14> cbl<7> in1<94> in2<94> sl<14> vdd vss wl<94> / cell_PIM
XI18084 bl<14> cbl<7> in1<95> in2<95> sl<14> vdd vss wl<95> / cell_PIM
XI18738 bl<14> cbl<7> in1<14> in2<14> sl<14> vdd vss wl<14> / cell_PIM
XI18737 bl<14> cbl<7> in1<10> in2<10> sl<14> vdd vss wl<10> / cell_PIM
XI17430 bl<6> cbl<3> in1<93> in2<93> sl<6> vdd vss wl<93> / cell_PIM
XI17429 bl<6> cbl<3> in1<94> in2<94> sl<6> vdd vss wl<94> / cell_PIM
XI18083 bl<14> cbl<7> in1<92> in2<92> sl<14> vdd vss wl<92> / cell_PIM
XI18731 bl<12> cbl<6> in1<14> in2<14> sl<12> vdd vss wl<14> / cell_PIM
XI18730 bl<12> cbl<6> in1<13> in2<13> sl<12> vdd vss wl<13> / cell_PIM
XI18729 bl<12> cbl<6> in1<12> in2<12> sl<12> vdd vss wl<12> / cell_PIM
XI18728 bl<12> cbl<6> in1<11> in2<11> sl<12> vdd vss wl<11> / cell_PIM
XI18727 bl<12> cbl<6> in1<10> in2<10> sl<12> vdd vss wl<10> / cell_PIM
XI18078 bl<12> cbl<6> in1<95> in2<95> sl<12> vdd vss wl<95> / cell_PIM
XI18077 bl<12> cbl<6> in1<94> in2<94> sl<12> vdd vss wl<94> / cell_PIM
XI18076 bl<12> cbl<6> in1<93> in2<93> sl<12> vdd vss wl<93> / cell_PIM
XI18075 bl<12> cbl<6> in1<92> in2<92> sl<12> vdd vss wl<92> / cell_PIM
XI17428 bl<6> cbl<3> in1<95> in2<95> sl<6> vdd vss wl<95> / cell_PIM
XI17427 bl<6> cbl<3> in1<92> in2<92> sl<6> vdd vss wl<92> / cell_PIM
XI17422 bl<4> cbl<2> in1<95> in2<95> sl<4> vdd vss wl<95> / cell_PIM
XI17421 bl<4> cbl<2> in1<94> in2<94> sl<4> vdd vss wl<94> / cell_PIM
XI17420 bl<4> cbl<2> in1<93> in2<93> sl<4> vdd vss wl<93> / cell_PIM
XI17419 bl<4> cbl<2> in1<92> in2<92> sl<4> vdd vss wl<92> / cell_PIM
XI18070 bl<10> cbl<5> in1<93> in2<93> sl<10> vdd vss wl<93> / cell_PIM
XI18069 bl<10> cbl<5> in1<94> in2<94> sl<10> vdd vss wl<94> / cell_PIM
XI18721 bl<10> cbl<5> in1<11> in2<11> sl<10> vdd vss wl<11> / cell_PIM
XI18720 bl<10> cbl<5> in1<12> in2<12> sl<10> vdd vss wl<12> / cell_PIM
XI18719 bl<10> cbl<5> in1<13> in2<13> sl<10> vdd vss wl<13> / cell_PIM
XI18068 bl<10> cbl<5> in1<95> in2<95> sl<10> vdd vss wl<95> / cell_PIM
XI18067 bl<10> cbl<5> in1<92> in2<92> sl<10> vdd vss wl<92> / cell_PIM
XI18718 bl<10> cbl<5> in1<14> in2<14> sl<10> vdd vss wl<14> / cell_PIM
XI18717 bl<10> cbl<5> in1<10> in2<10> sl<10> vdd vss wl<10> / cell_PIM
XI17413 bl<6> cbl<3> in1<97> in2<97> sl<6> vdd vss wl<97> / cell_PIM
XI17412 bl<6> cbl<3> in1<98> in2<98> sl<6> vdd vss wl<98> / cell_PIM
XI17411 bl<6> cbl<3> in1<99> in2<99> sl<6> vdd vss wl<99> / cell_PIM
XI17410 bl<6> cbl<3> in1<100> in2<100> sl<6> vdd vss wl<100> / cell_PIM
XI17409 bl<6> cbl<3> in1<96> in2<96> sl<6> vdd vss wl<96> / cell_PIM
XI18062 bl<8> cbl<4> in1<95> in2<95> sl<8> vdd vss wl<95> / cell_PIM
XI18061 bl<8> cbl<4> in1<94> in2<94> sl<8> vdd vss wl<94> / cell_PIM
XI18060 bl<8> cbl<4> in1<93> in2<93> sl<8> vdd vss wl<93> / cell_PIM
XI18059 bl<8> cbl<4> in1<92> in2<92> sl<8> vdd vss wl<92> / cell_PIM
XI18711 bl<8> cbl<4> in1<14> in2<14> sl<8> vdd vss wl<14> / cell_PIM
XI18710 bl<8> cbl<4> in1<13> in2<13> sl<8> vdd vss wl<13> / cell_PIM
XI18709 bl<8> cbl<4> in1<12> in2<12> sl<8> vdd vss wl<12> / cell_PIM
XI18708 bl<8> cbl<4> in1<11> in2<11> sl<8> vdd vss wl<11> / cell_PIM
XI18707 bl<8> cbl<4> in1<10> in2<10> sl<8> vdd vss wl<10> / cell_PIM
XI17403 bl<4> cbl<2> in1<100> in2<100> sl<4> vdd vss wl<100> / cell_PIM
XI17402 bl<4> cbl<2> in1<99> in2<99> sl<4> vdd vss wl<99> / cell_PIM
XI17401 bl<4> cbl<2> in1<98> in2<98> sl<4> vdd vss wl<98> / cell_PIM
XI17400 bl<4> cbl<2> in1<97> in2<97> sl<4> vdd vss wl<97> / cell_PIM
XI17399 bl<4> cbl<2> in1<96> in2<96> sl<4> vdd vss wl<96> / cell_PIM
XI18053 bl<14> cbl<7> in1<97> in2<97> sl<14> vdd vss wl<97> / cell_PIM
XI18052 bl<14> cbl<7> in1<98> in2<98> sl<14> vdd vss wl<98> / cell_PIM
XI18051 bl<14> cbl<7> in1<99> in2<99> sl<14> vdd vss wl<99> / cell_PIM
XI18050 bl<14> cbl<7> in1<100> in2<100> sl<14> vdd vss wl<100> / cell_PIM
XI18049 bl<14> cbl<7> in1<96> in2<96> sl<14> vdd vss wl<96> / cell_PIM
XI18701 bl<14> cbl<7> in1<16> in2<16> sl<14> vdd vss wl<16> / cell_PIM
XI18700 bl<14> cbl<7> in1<17> in2<17> sl<14> vdd vss wl<17> / cell_PIM
XI18699 bl<14> cbl<7> in1<18> in2<18> sl<14> vdd vss wl<18> / cell_PIM
XI18698 bl<14> cbl<7> in1<19> in2<19> sl<14> vdd vss wl<19> / cell_PIM
XI18697 bl<14> cbl<7> in1<15> in2<15> sl<14> vdd vss wl<15> / cell_PIM
XI17393 bl<6> cbl<3> in1<102> in2<102> sl<6> vdd vss wl<102> / cell_PIM
XI17392 bl<6> cbl<3> in1<103> in2<103> sl<6> vdd vss wl<103> / cell_PIM
XI17391 bl<6> cbl<3> in1<104> in2<104> sl<6> vdd vss wl<104> / cell_PIM
XI17390 bl<6> cbl<3> in1<105> in2<105> sl<6> vdd vss wl<105> / cell_PIM
XI17389 bl<6> cbl<3> in1<101> in2<101> sl<6> vdd vss wl<101> / cell_PIM
XI18043 bl<12> cbl<6> in1<100> in2<100> sl<12> vdd vss wl<100> / cell_PIM
XI18042 bl<12> cbl<6> in1<99> in2<99> sl<12> vdd vss wl<99> / cell_PIM
XI18041 bl<12> cbl<6> in1<98> in2<98> sl<12> vdd vss wl<98> / cell_PIM
XI18040 bl<12> cbl<6> in1<97> in2<97> sl<12> vdd vss wl<97> / cell_PIM
XI18039 bl<12> cbl<6> in1<96> in2<96> sl<12> vdd vss wl<96> / cell_PIM
XI18691 bl<12> cbl<6> in1<19> in2<19> sl<12> vdd vss wl<19> / cell_PIM
XI18690 bl<12> cbl<6> in1<18> in2<18> sl<12> vdd vss wl<18> / cell_PIM
XI18689 bl<12> cbl<6> in1<17> in2<17> sl<12> vdd vss wl<17> / cell_PIM
XI18688 bl<12> cbl<6> in1<16> in2<16> sl<12> vdd vss wl<16> / cell_PIM
XI18687 bl<12> cbl<6> in1<15> in2<15> sl<12> vdd vss wl<15> / cell_PIM
XI17383 bl<4> cbl<2> in1<105> in2<105> sl<4> vdd vss wl<105> / cell_PIM
XI17382 bl<4> cbl<2> in1<104> in2<104> sl<4> vdd vss wl<104> / cell_PIM
XI17381 bl<4> cbl<2> in1<103> in2<103> sl<4> vdd vss wl<103> / cell_PIM
XI17380 bl<4> cbl<2> in1<102> in2<102> sl<4> vdd vss wl<102> / cell_PIM
XI17379 bl<4> cbl<2> in1<101> in2<101> sl<4> vdd vss wl<101> / cell_PIM
XI18033 bl<10> cbl<5> in1<97> in2<97> sl<10> vdd vss wl<97> / cell_PIM
XI18032 bl<10> cbl<5> in1<98> in2<98> sl<10> vdd vss wl<98> / cell_PIM
XI18031 bl<10> cbl<5> in1<99> in2<99> sl<10> vdd vss wl<99> / cell_PIM
XI18030 bl<10> cbl<5> in1<100> in2<100> sl<10> vdd vss wl<100> / cell_PIM
XI18029 bl<10> cbl<5> in1<96> in2<96> sl<10> vdd vss wl<96> / cell_PIM
XI18681 bl<10> cbl<5> in1<16> in2<16> sl<10> vdd vss wl<16> / cell_PIM
XI18680 bl<10> cbl<5> in1<17> in2<17> sl<10> vdd vss wl<17> / cell_PIM
XI18679 bl<10> cbl<5> in1<18> in2<18> sl<10> vdd vss wl<18> / cell_PIM
XI18678 bl<10> cbl<5> in1<19> in2<19> sl<10> vdd vss wl<19> / cell_PIM
XI18677 bl<10> cbl<5> in1<15> in2<15> sl<10> vdd vss wl<15> / cell_PIM
XI17373 bl<6> cbl<3> in1<107> in2<107> sl<6> vdd vss wl<107> / cell_PIM
XI17372 bl<6> cbl<3> in1<108> in2<108> sl<6> vdd vss wl<108> / cell_PIM
XI17371 bl<6> cbl<3> in1<109> in2<109> sl<6> vdd vss wl<109> / cell_PIM
XI17370 bl<6> cbl<3> in1<110> in2<110> sl<6> vdd vss wl<110> / cell_PIM
XI17369 bl<6> cbl<3> in1<106> in2<106> sl<6> vdd vss wl<106> / cell_PIM
XI18023 bl<8> cbl<4> in1<100> in2<100> sl<8> vdd vss wl<100> / cell_PIM
XI18022 bl<8> cbl<4> in1<99> in2<99> sl<8> vdd vss wl<99> / cell_PIM
XI18021 bl<8> cbl<4> in1<98> in2<98> sl<8> vdd vss wl<98> / cell_PIM
XI18020 bl<8> cbl<4> in1<97> in2<97> sl<8> vdd vss wl<97> / cell_PIM
XI18019 bl<8> cbl<4> in1<96> in2<96> sl<8> vdd vss wl<96> / cell_PIM
XI18671 bl<8> cbl<4> in1<19> in2<19> sl<8> vdd vss wl<19> / cell_PIM
XI18670 bl<8> cbl<4> in1<18> in2<18> sl<8> vdd vss wl<18> / cell_PIM
XI18669 bl<8> cbl<4> in1<17> in2<17> sl<8> vdd vss wl<17> / cell_PIM
XI18668 bl<8> cbl<4> in1<16> in2<16> sl<8> vdd vss wl<16> / cell_PIM
XI18667 bl<8> cbl<4> in1<15> in2<15> sl<8> vdd vss wl<15> / cell_PIM
XI17363 bl<4> cbl<2> in1<110> in2<110> sl<4> vdd vss wl<110> / cell_PIM
XI17362 bl<4> cbl<2> in1<109> in2<109> sl<4> vdd vss wl<109> / cell_PIM
XI17361 bl<4> cbl<2> in1<108> in2<108> sl<4> vdd vss wl<108> / cell_PIM
XI17360 bl<4> cbl<2> in1<107> in2<107> sl<4> vdd vss wl<107> / cell_PIM
XI17359 bl<4> cbl<2> in1<106> in2<106> sl<4> vdd vss wl<106> / cell_PIM
XI18013 bl<14> cbl<7> in1<102> in2<102> sl<14> vdd vss wl<102> / cell_PIM
XI18012 bl<14> cbl<7> in1<103> in2<103> sl<14> vdd vss wl<103> / cell_PIM
XI18011 bl<14> cbl<7> in1<104> in2<104> sl<14> vdd vss wl<104> / cell_PIM
XI18010 bl<14> cbl<7> in1<105> in2<105> sl<14> vdd vss wl<105> / cell_PIM
XI18009 bl<14> cbl<7> in1<101> in2<101> sl<14> vdd vss wl<101> / cell_PIM
XI18661 bl<14> cbl<7> in1<21> in2<21> sl<14> vdd vss wl<21> / cell_PIM
XI18660 bl<14> cbl<7> in1<22> in2<22> sl<14> vdd vss wl<22> / cell_PIM
XI18659 bl<14> cbl<7> in1<23> in2<23> sl<14> vdd vss wl<23> / cell_PIM
XI18658 bl<14> cbl<7> in1<24> in2<24> sl<14> vdd vss wl<24> / cell_PIM
XI18657 bl<14> cbl<7> in1<20> in2<20> sl<14> vdd vss wl<20> / cell_PIM
XI17353 bl<6> cbl<3> in1<112> in2<112> sl<6> vdd vss wl<112> / cell_PIM
XI17352 bl<6> cbl<3> in1<113> in2<113> sl<6> vdd vss wl<113> / cell_PIM
XI17351 bl<6> cbl<3> in1<114> in2<114> sl<6> vdd vss wl<114> / cell_PIM
XI17350 bl<6> cbl<3> in1<115> in2<115> sl<6> vdd vss wl<115> / cell_PIM
XI17349 bl<6> cbl<3> in1<111> in2<111> sl<6> vdd vss wl<111> / cell_PIM
XI18003 bl<12> cbl<6> in1<105> in2<105> sl<12> vdd vss wl<105> / cell_PIM
XI18002 bl<12> cbl<6> in1<104> in2<104> sl<12> vdd vss wl<104> / cell_PIM
XI18001 bl<12> cbl<6> in1<103> in2<103> sl<12> vdd vss wl<103> / cell_PIM
XI18000 bl<12> cbl<6> in1<102> in2<102> sl<12> vdd vss wl<102> / cell_PIM
XI17999 bl<12> cbl<6> in1<101> in2<101> sl<12> vdd vss wl<101> / cell_PIM
XI18651 bl<12> cbl<6> in1<24> in2<24> sl<12> vdd vss wl<24> / cell_PIM
XI18650 bl<12> cbl<6> in1<23> in2<23> sl<12> vdd vss wl<23> / cell_PIM
XI18649 bl<12> cbl<6> in1<22> in2<22> sl<12> vdd vss wl<22> / cell_PIM
XI18648 bl<12> cbl<6> in1<21> in2<21> sl<12> vdd vss wl<21> / cell_PIM
XI18647 bl<12> cbl<6> in1<20> in2<20> sl<12> vdd vss wl<20> / cell_PIM
XI17343 bl<4> cbl<2> in1<115> in2<115> sl<4> vdd vss wl<115> / cell_PIM
XI17342 bl<4> cbl<2> in1<114> in2<114> sl<4> vdd vss wl<114> / cell_PIM
XI17341 bl<4> cbl<2> in1<113> in2<113> sl<4> vdd vss wl<113> / cell_PIM
XI17340 bl<4> cbl<2> in1<112> in2<112> sl<4> vdd vss wl<112> / cell_PIM
XI17339 bl<4> cbl<2> in1<111> in2<111> sl<4> vdd vss wl<111> / cell_PIM
XI17993 bl<10> cbl<5> in1<102> in2<102> sl<10> vdd vss wl<102> / cell_PIM
XI17992 bl<10> cbl<5> in1<103> in2<103> sl<10> vdd vss wl<103> / cell_PIM
XI17991 bl<10> cbl<5> in1<104> in2<104> sl<10> vdd vss wl<104> / cell_PIM
XI17990 bl<10> cbl<5> in1<105> in2<105> sl<10> vdd vss wl<105> / cell_PIM
XI17989 bl<10> cbl<5> in1<101> in2<101> sl<10> vdd vss wl<101> / cell_PIM
XI18641 bl<10> cbl<5> in1<21> in2<21> sl<10> vdd vss wl<21> / cell_PIM
XI18640 bl<10> cbl<5> in1<22> in2<22> sl<10> vdd vss wl<22> / cell_PIM
XI18639 bl<10> cbl<5> in1<23> in2<23> sl<10> vdd vss wl<23> / cell_PIM
XI17334 bl<6> cbl<3> in1<117> in2<117> sl<6> vdd vss wl<117> / cell_PIM
XI18638 bl<10> cbl<5> in1<24> in2<24> sl<10> vdd vss wl<24> / cell_PIM
XI18637 bl<10> cbl<5> in1<20> in2<20> sl<10> vdd vss wl<20> / cell_PIM
XI16874 bl<0> cbl<0> in1<95> in2<95> sl<0> vdd vss wl<95> / cell_PIM
XI16873 bl<0> cbl<0> in1<94> in2<94> sl<0> vdd vss wl<94> / cell_PIM
XI16871 bl<0> cbl<0> in1<92> in2<92> sl<0> vdd vss wl<92> / cell_PIM
XI16870 bl<0> cbl<0> in1<91> in2<91> sl<0> vdd vss wl<91> / cell_PIM
XI16868 bl<0> cbl<0> in1<89> in2<89> sl<0> vdd vss wl<89> / cell_PIM
XI16867 bl<0> cbl<0> in1<88> in2<88> sl<0> vdd vss wl<88> / cell_PIM
XI16865 bl<0> cbl<0> in1<86> in2<86> sl<0> vdd vss wl<86> / cell_PIM
XI16864 bl<0> cbl<0> in1<85> in2<85> sl<0> vdd vss wl<85> / cell_PIM
XI16862 bl<0> cbl<0> in1<83> in2<83> sl<0> vdd vss wl<83> / cell_PIM
XI16861 bl<0> cbl<0> in1<82> in2<82> sl<0> vdd vss wl<82> / cell_PIM
XI16859 bl<0> cbl<0> in1<80> in2<80> sl<0> vdd vss wl<80> / cell_PIM
XI16858 bl<0> cbl<0> in1<79> in2<79> sl<0> vdd vss wl<79> / cell_PIM
XI16856 bl<0> cbl<0> in1<77> in2<77> sl<0> vdd vss wl<77> / cell_PIM
XI16855 bl<0> cbl<0> in1<76> in2<76> sl<0> vdd vss wl<76> / cell_PIM
XI16853 bl<0> cbl<0> in1<74> in2<74> sl<0> vdd vss wl<74> / cell_PIM
XI16852 bl<0> cbl<0> in1<73> in2<73> sl<0> vdd vss wl<73> / cell_PIM
XI16850 bl<0> cbl<0> in1<71> in2<71> sl<0> vdd vss wl<71> / cell_PIM
XI16849 bl<0> cbl<0> in1<70> in2<70> sl<0> vdd vss wl<70> / cell_PIM
XI16812 bl<0> cbl<0> in1<33> in2<33> sl<0> vdd vss wl<33> / cell_PIM
XI16811 bl<0> cbl<0> in1<32> in2<32> sl<0> vdd vss wl<32> / cell_PIM
XI16809 bl<0> cbl<0> in1<30> in2<30> sl<0> vdd vss wl<30> / cell_PIM
XI16808 bl<0> cbl<0> in1<29> in2<29> sl<0> vdd vss wl<29> / cell_PIM
XI16806 bl<0> cbl<0> in1<27> in2<27> sl<0> vdd vss wl<27> / cell_PIM
XI16805 bl<0> cbl<0> in1<26> in2<26> sl<0> vdd vss wl<26> / cell_PIM
XI16803 bl<0> cbl<0> in1<24> in2<24> sl<0> vdd vss wl<24> / cell_PIM
XI16802 bl<0> cbl<0> in1<23> in2<23> sl<0> vdd vss wl<23> / cell_PIM
XI16800 bl<0> cbl<0> in1<21> in2<21> sl<0> vdd vss wl<21> / cell_PIM
XI16799 bl<0> cbl<0> in1<20> in2<20> sl<0> vdd vss wl<20> / cell_PIM
XI16797 bl<0> cbl<0> in1<18> in2<18> sl<0> vdd vss wl<18> / cell_PIM
XI16796 bl<0> cbl<0> in1<17> in2<17> sl<0> vdd vss wl<17> / cell_PIM
XI16794 bl<0> cbl<0> in1<15> in2<15> sl<0> vdd vss wl<15> / cell_PIM
XI16793 bl<0> cbl<0> in1<14> in2<14> sl<0> vdd vss wl<14> / cell_PIM
XI24869 bl<62> cbl<31> in1<3> in2<3> sl<62> vdd vss wl<3> / cell_PIM
XI24868 bl<62> cbl<31> in1<4> in2<4> sl<62> vdd vss wl<4> / cell_PIM
XI24867 bl<62> cbl<31> in1<6> in2<6> sl<62> vdd vss wl<6> / cell_PIM
XI24866 bl<62> cbl<31> in1<7> in2<7> sl<62> vdd vss wl<7> / cell_PIM
XI24865 bl<62> cbl<31> in1<5> in2<5> sl<62> vdd vss wl<5> / cell_PIM
XI24218 bl<54> cbl<27> in1<26> in2<26> sl<54> vdd vss wl<26> / cell_PIM
XI24859 bl<60> cbl<30> in1<4> in2<4> sl<60> vdd vss wl<4> / cell_PIM
XI24208 bl<52> cbl<26> in1<26> in2<26> sl<52> vdd vss wl<26> / cell_PIM
XI24857 bl<60> cbl<30> in1<7> in2<7> sl<60> vdd vss wl<7> / cell_PIM
XI24856 bl<60> cbl<30> in1<6> in2<6> sl<60> vdd vss wl<6> / cell_PIM
XI24855 bl<60> cbl<30> in1<5> in2<5> sl<60> vdd vss wl<5> / cell_PIM
XI24858 bl<60> cbl<30> in1<3> in2<3> sl<60> vdd vss wl<3> / cell_PIM
XI24849 bl<58> cbl<29> in1<3> in2<3> sl<58> vdd vss wl<3> / cell_PIM
XI24848 bl<58> cbl<29> in1<4> in2<4> sl<58> vdd vss wl<4> / cell_PIM
XI24847 bl<58> cbl<29> in1<6> in2<6> sl<58> vdd vss wl<6> / cell_PIM
XI24846 bl<58> cbl<29> in1<7> in2<7> sl<58> vdd vss wl<7> / cell_PIM
XI24845 bl<58> cbl<29> in1<5> in2<5> sl<58> vdd vss wl<5> / cell_PIM
XI24198 bl<50> cbl<25> in1<26> in2<26> sl<50> vdd vss wl<26> / cell_PIM
XI24839 bl<56> cbl<28> in1<3> in2<3> sl<56> vdd vss wl<3> / cell_PIM
XI24188 bl<48> cbl<24> in1<26> in2<26> sl<48> vdd vss wl<26> / cell_PIM
XI24837 bl<56> cbl<28> in1<6> in2<6> sl<56> vdd vss wl<6> / cell_PIM
XI24836 bl<56> cbl<28> in1<7> in2<7> sl<56> vdd vss wl<7> / cell_PIM
XI24835 bl<56> cbl<28> in1<5> in2<5> sl<56> vdd vss wl<5> / cell_PIM
XI24838 bl<56> cbl<28> in1<4> in2<4> sl<56> vdd vss wl<4> / cell_PIM
XI24829 bl<54> cbl<27> in1<3> in2<3> sl<54> vdd vss wl<3> / cell_PIM
XI24828 bl<54> cbl<27> in1<4> in2<4> sl<54> vdd vss wl<4> / cell_PIM
XI24827 bl<54> cbl<27> in1<6> in2<6> sl<54> vdd vss wl<6> / cell_PIM
XI24826 bl<54> cbl<27> in1<7> in2<7> sl<54> vdd vss wl<7> / cell_PIM
XI24825 bl<54> cbl<27> in1<5> in2<5> sl<54> vdd vss wl<5> / cell_PIM
XI24178 bl<46> cbl<23> in1<26> in2<26> sl<46> vdd vss wl<26> / cell_PIM
XI24819 bl<52> cbl<26> in1<4> in2<4> sl<52> vdd vss wl<4> / cell_PIM
XI24168 bl<44> cbl<22> in1<26> in2<26> sl<44> vdd vss wl<26> / cell_PIM
XI24817 bl<52> cbl<26> in1<7> in2<7> sl<52> vdd vss wl<7> / cell_PIM
XI24816 bl<52> cbl<26> in1<6> in2<6> sl<52> vdd vss wl<6> / cell_PIM
XI24815 bl<52> cbl<26> in1<5> in2<5> sl<52> vdd vss wl<5> / cell_PIM
XI24818 bl<52> cbl<26> in1<3> in2<3> sl<52> vdd vss wl<3> / cell_PIM
XI24809 bl<50> cbl<25> in1<3> in2<3> sl<50> vdd vss wl<3> / cell_PIM
XI24808 bl<50> cbl<25> in1<4> in2<4> sl<50> vdd vss wl<4> / cell_PIM
XI24807 bl<50> cbl<25> in1<6> in2<6> sl<50> vdd vss wl<6> / cell_PIM
XI24806 bl<50> cbl<25> in1<7> in2<7> sl<50> vdd vss wl<7> / cell_PIM
XI24805 bl<50> cbl<25> in1<5> in2<5> sl<50> vdd vss wl<5> / cell_PIM
XI24158 bl<42> cbl<21> in1<26> in2<26> sl<42> vdd vss wl<26> / cell_PIM
XI24799 bl<48> cbl<24> in1<4> in2<4> sl<48> vdd vss wl<4> / cell_PIM
XI24148 bl<40> cbl<20> in1<26> in2<26> sl<40> vdd vss wl<26> / cell_PIM
XI24797 bl<48> cbl<24> in1<7> in2<7> sl<48> vdd vss wl<7> / cell_PIM
XI24796 bl<48> cbl<24> in1<6> in2<6> sl<48> vdd vss wl<6> / cell_PIM
XI24795 bl<48> cbl<24> in1<5> in2<5> sl<48> vdd vss wl<5> / cell_PIM
XI24798 bl<48> cbl<24> in1<3> in2<3> sl<48> vdd vss wl<3> / cell_PIM
XI22403 bl<62> cbl<31> in1<82> in2<82> sl<62> vdd vss wl<82> / cell_PIM
XI23020 bl<32> cbl<16> in1<59> in2<59> sl<32> vdd vss wl<59> / cell_PIM
XI23019 bl<32> cbl<16> in1<58> in2<58> sl<32> vdd vss wl<58> / cell_PIM
XI23573 bl<46> cbl<23> in1<41> in2<41> sl<46> vdd vss wl<41> / cell_PIM
XI23572 bl<46> cbl<23> in1<42> in2<42> sl<46> vdd vss wl<42> / cell_PIM
XI23571 bl<46> cbl<23> in1<43> in2<43> sl<46> vdd vss wl<43> / cell_PIM
XI23570 bl<46> cbl<23> in1<45> in2<45> sl<46> vdd vss wl<45> / cell_PIM
XI23569 bl<46> cbl<23> in1<44> in2<44> sl<46> vdd vss wl<44> / cell_PIM
XI24221 bl<54> cbl<27> in1<22> in2<22> sl<54> vdd vss wl<22> / cell_PIM
XI24220 bl<54> cbl<27> in1<23> in2<23> sl<54> vdd vss wl<23> / cell_PIM
XI24219 bl<54> cbl<27> in1<24> in2<24> sl<54> vdd vss wl<24> / cell_PIM
XI24217 bl<54> cbl<27> in1<25> in2<25> sl<54> vdd vss wl<25> / cell_PIM
XI23014 bl<62> cbl<31> in1<61> in2<61> sl<62> vdd vss wl<61> / cell_PIM
XI23013 bl<62> cbl<31> in1<62> in2<62> sl<62> vdd vss wl<62> / cell_PIM
XI22398 bl<60> cbl<30> in1<81> in2<81> sl<60> vdd vss wl<81> / cell_PIM
XI23012 bl<62> cbl<31> in1<64> in2<64> sl<62> vdd vss wl<64> / cell_PIM
XI23011 bl<62> cbl<31> in1<63> in2<63> sl<62> vdd vss wl<63> / cell_PIM
XI23563 bl<44> cbl<22> in1<43> in2<43> sl<44> vdd vss wl<43> / cell_PIM
XI23562 bl<44> cbl<22> in1<42> in2<42> sl<44> vdd vss wl<42> / cell_PIM
XI23561 bl<44> cbl<22> in1<41> in2<41> sl<44> vdd vss wl<41> / cell_PIM
XI23560 bl<44> cbl<22> in1<45> in2<45> sl<44> vdd vss wl<45> / cell_PIM
XI23559 bl<44> cbl<22> in1<44> in2<44> sl<44> vdd vss wl<44> / cell_PIM
XI24211 bl<52> cbl<26> in1<24> in2<24> sl<52> vdd vss wl<24> / cell_PIM
XI24210 bl<52> cbl<26> in1<23> in2<23> sl<52> vdd vss wl<23> / cell_PIM
XI24209 bl<52> cbl<26> in1<22> in2<22> sl<52> vdd vss wl<22> / cell_PIM
XI22388 bl<58> cbl<29> in1<83> in2<83> sl<58> vdd vss wl<83> / cell_PIM
XI23006 bl<60> cbl<30> in1<62> in2<62> sl<60> vdd vss wl<62> / cell_PIM
XI23005 bl<60> cbl<30> in1<61> in2<61> sl<60> vdd vss wl<61> / cell_PIM
XI24207 bl<52> cbl<26> in1<25> in2<25> sl<52> vdd vss wl<25> / cell_PIM
XI23004 bl<60> cbl<30> in1<64> in2<64> sl<60> vdd vss wl<64> / cell_PIM
XI23003 bl<60> cbl<30> in1<63> in2<63> sl<60> vdd vss wl<63> / cell_PIM
XI23553 bl<42> cbl<21> in1<41> in2<41> sl<42> vdd vss wl<41> / cell_PIM
XI23552 bl<42> cbl<21> in1<42> in2<42> sl<42> vdd vss wl<42> / cell_PIM
XI23551 bl<42> cbl<21> in1<43> in2<43> sl<42> vdd vss wl<43> / cell_PIM
XI23550 bl<42> cbl<21> in1<45> in2<45> sl<42> vdd vss wl<45> / cell_PIM
XI23549 bl<42> cbl<21> in1<44> in2<44> sl<42> vdd vss wl<44> / cell_PIM
XI24201 bl<50> cbl<25> in1<22> in2<22> sl<50> vdd vss wl<22> / cell_PIM
XI24200 bl<50> cbl<25> in1<23> in2<23> sl<50> vdd vss wl<23> / cell_PIM
XI24199 bl<50> cbl<25> in1<24> in2<24> sl<50> vdd vss wl<24> / cell_PIM
XI24197 bl<50> cbl<25> in1<25> in2<25> sl<50> vdd vss wl<25> / cell_PIM
XI22998 bl<58> cbl<29> in1<61> in2<61> sl<58> vdd vss wl<61> / cell_PIM
XI22997 bl<58> cbl<29> in1<62> in2<62> sl<58> vdd vss wl<62> / cell_PIM
XI22373 bl<54> cbl<27> in1<81> in2<81> sl<54> vdd vss wl<81> / cell_PIM
XI22996 bl<58> cbl<29> in1<64> in2<64> sl<58> vdd vss wl<64> / cell_PIM
XI22995 bl<58> cbl<29> in1<63> in2<63> sl<58> vdd vss wl<63> / cell_PIM
XI23543 bl<40> cbl<20> in1<41> in2<41> sl<40> vdd vss wl<41> / cell_PIM
XI23542 bl<40> cbl<20> in1<42> in2<42> sl<40> vdd vss wl<42> / cell_PIM
XI23541 bl<40> cbl<20> in1<43> in2<43> sl<40> vdd vss wl<43> / cell_PIM
XI23540 bl<40> cbl<20> in1<45> in2<45> sl<40> vdd vss wl<45> / cell_PIM
XI23539 bl<40> cbl<20> in1<44> in2<44> sl<40> vdd vss wl<44> / cell_PIM
XI24191 bl<48> cbl<24> in1<24> in2<24> sl<48> vdd vss wl<24> / cell_PIM
XI24190 bl<48> cbl<24> in1<23> in2<23> sl<48> vdd vss wl<23> / cell_PIM
XI24189 bl<48> cbl<24> in1<22> in2<22> sl<48> vdd vss wl<22> / cell_PIM
XI22990 bl<56> cbl<28> in1<61> in2<61> sl<56> vdd vss wl<61> / cell_PIM
XI22989 bl<56> cbl<28> in1<62> in2<62> sl<56> vdd vss wl<62> / cell_PIM
XI24187 bl<48> cbl<24> in1<25> in2<25> sl<48> vdd vss wl<25> / cell_PIM
XI22363 bl<52> cbl<26> in1<82> in2<82> sl<52> vdd vss wl<82> / cell_PIM
XI22988 bl<56> cbl<28> in1<64> in2<64> sl<56> vdd vss wl<64> / cell_PIM
XI22987 bl<56> cbl<28> in1<63> in2<63> sl<56> vdd vss wl<63> / cell_PIM
XI23533 bl<38> cbl<19> in1<41> in2<41> sl<38> vdd vss wl<41> / cell_PIM
XI23532 bl<38> cbl<19> in1<42> in2<42> sl<38> vdd vss wl<42> / cell_PIM
XI23531 bl<38> cbl<19> in1<43> in2<43> sl<38> vdd vss wl<43> / cell_PIM
XI23530 bl<38> cbl<19> in1<45> in2<45> sl<38> vdd vss wl<45> / cell_PIM
XI23529 bl<38> cbl<19> in1<44> in2<44> sl<38> vdd vss wl<44> / cell_PIM
XI24181 bl<46> cbl<23> in1<22> in2<22> sl<46> vdd vss wl<22> / cell_PIM
XI24180 bl<46> cbl<23> in1<23> in2<23> sl<46> vdd vss wl<23> / cell_PIM
XI24179 bl<46> cbl<23> in1<24> in2<24> sl<46> vdd vss wl<24> / cell_PIM
XI24177 bl<46> cbl<23> in1<25> in2<25> sl<46> vdd vss wl<25> / cell_PIM
XI22982 bl<54> cbl<27> in1<61> in2<61> sl<54> vdd vss wl<61> / cell_PIM
XI22981 bl<54> cbl<27> in1<62> in2<62> sl<54> vdd vss wl<62> / cell_PIM
XI22358 bl<50> cbl<25> in1<80> in2<80> sl<50> vdd vss wl<80> / cell_PIM
XI22980 bl<54> cbl<27> in1<64> in2<64> sl<54> vdd vss wl<64> / cell_PIM
XI22979 bl<54> cbl<27> in1<63> in2<63> sl<54> vdd vss wl<63> / cell_PIM
XI23523 bl<36> cbl<18> in1<43> in2<43> sl<36> vdd vss wl<43> / cell_PIM
XI23522 bl<36> cbl<18> in1<42> in2<42> sl<36> vdd vss wl<42> / cell_PIM
XI23521 bl<36> cbl<18> in1<41> in2<41> sl<36> vdd vss wl<41> / cell_PIM
XI23520 bl<36> cbl<18> in1<45> in2<45> sl<36> vdd vss wl<45> / cell_PIM
XI23519 bl<36> cbl<18> in1<44> in2<44> sl<36> vdd vss wl<44> / cell_PIM
XI24171 bl<44> cbl<22> in1<24> in2<24> sl<44> vdd vss wl<24> / cell_PIM
XI24170 bl<44> cbl<22> in1<23> in2<23> sl<44> vdd vss wl<23> / cell_PIM
XI24169 bl<44> cbl<22> in1<22> in2<22> sl<44> vdd vss wl<22> / cell_PIM
XI22348 bl<48> cbl<24> in1<83> in2<83> sl<48> vdd vss wl<83> / cell_PIM
XI22974 bl<52> cbl<26> in1<62> in2<62> sl<52> vdd vss wl<62> / cell_PIM
XI22973 bl<52> cbl<26> in1<61> in2<61> sl<52> vdd vss wl<61> / cell_PIM
XI24167 bl<44> cbl<22> in1<25> in2<25> sl<44> vdd vss wl<25> / cell_PIM
XI22972 bl<52> cbl<26> in1<64> in2<64> sl<52> vdd vss wl<64> / cell_PIM
XI22971 bl<52> cbl<26> in1<63> in2<63> sl<52> vdd vss wl<63> / cell_PIM
XI23513 bl<34> cbl<17> in1<41> in2<41> sl<34> vdd vss wl<41> / cell_PIM
XI23512 bl<34> cbl<17> in1<42> in2<42> sl<34> vdd vss wl<42> / cell_PIM
XI23511 bl<34> cbl<17> in1<43> in2<43> sl<34> vdd vss wl<43> / cell_PIM
XI23510 bl<34> cbl<17> in1<45> in2<45> sl<34> vdd vss wl<45> / cell_PIM
XI23509 bl<34> cbl<17> in1<44> in2<44> sl<34> vdd vss wl<44> / cell_PIM
XI24161 bl<42> cbl<21> in1<22> in2<22> sl<42> vdd vss wl<22> / cell_PIM
XI24160 bl<42> cbl<21> in1<23> in2<23> sl<42> vdd vss wl<23> / cell_PIM
XI24159 bl<42> cbl<21> in1<24> in2<24> sl<42> vdd vss wl<24> / cell_PIM
XI24157 bl<42> cbl<21> in1<25> in2<25> sl<42> vdd vss wl<25> / cell_PIM
XI22966 bl<50> cbl<25> in1<61> in2<61> sl<50> vdd vss wl<61> / cell_PIM
XI22965 bl<50> cbl<25> in1<62> in2<62> sl<50> vdd vss wl<62> / cell_PIM
XI22333 bl<44> cbl<22> in1<80> in2<80> sl<44> vdd vss wl<80> / cell_PIM
XI22964 bl<50> cbl<25> in1<64> in2<64> sl<50> vdd vss wl<64> / cell_PIM
XI22963 bl<50> cbl<25> in1<63> in2<63> sl<50> vdd vss wl<63> / cell_PIM
XI23503 bl<32> cbl<16> in1<43> in2<43> sl<32> vdd vss wl<43> / cell_PIM
XI23502 bl<32> cbl<16> in1<42> in2<42> sl<32> vdd vss wl<42> / cell_PIM
XI23501 bl<32> cbl<16> in1<41> in2<41> sl<32> vdd vss wl<41> / cell_PIM
XI23500 bl<32> cbl<16> in1<45> in2<45> sl<32> vdd vss wl<45> / cell_PIM
XI23499 bl<32> cbl<16> in1<44> in2<44> sl<32> vdd vss wl<44> / cell_PIM
XI24151 bl<40> cbl<20> in1<22> in2<22> sl<40> vdd vss wl<22> / cell_PIM
XI24150 bl<40> cbl<20> in1<23> in2<23> sl<40> vdd vss wl<23> / cell_PIM
XI24149 bl<40> cbl<20> in1<24> in2<24> sl<40> vdd vss wl<24> / cell_PIM
XI22958 bl<48> cbl<24> in1<62> in2<62> sl<48> vdd vss wl<62> / cell_PIM
XI22957 bl<48> cbl<24> in1<61> in2<61> sl<48> vdd vss wl<61> / cell_PIM
XI24147 bl<40> cbl<20> in1<25> in2<25> sl<40> vdd vss wl<25> / cell_PIM
XI21099 bl<44> cbl<22> in1<119> in2<119> sl<44> vdd vss wl<119> / cell_PIM
XI21753 bl<54> cbl<27> in1<101> in2<101> sl<54> vdd vss wl<101> / cell_PIM
XI22397 bl<60> cbl<30> in1<80> in2<80> sl<60> vdd vss wl<80> / cell_PIM
XI22396 bl<60> cbl<30> in1<83> in2<83> sl<60> vdd vss wl<83> / cell_PIM
XI22395 bl<60> cbl<30> in1<82> in2<82> sl<60> vdd vss wl<82> / cell_PIM
XI21747 bl<52> cbl<26> in1<100> in2<100> sl<52> vdd vss wl<100> / cell_PIM
XI21746 bl<52> cbl<26> in1<99> in2<99> sl<52> vdd vss wl<99> / cell_PIM
XI21745 bl<52> cbl<26> in1<103> in2<103> sl<52> vdd vss wl<103> / cell_PIM
XI21744 bl<52> cbl<26> in1<102> in2<102> sl<52> vdd vss wl<102> / cell_PIM
XI21098 bl<44> cbl<22> in1<118> in2<118> sl<44> vdd vss wl<118> / cell_PIM
XI21097 bl<44> cbl<22> in1<122> in2<122> sl<44> vdd vss wl<122> / cell_PIM
XI21096 bl<44> cbl<22> in1<121> in2<121> sl<44> vdd vss wl<121> / cell_PIM
XI21095 bl<44> cbl<22> in1<120> in2<120> sl<44> vdd vss wl<120> / cell_PIM
XI21089 bl<42> cbl<21> in1<118> in2<118> sl<42> vdd vss wl<118> / cell_PIM
XI21743 bl<52> cbl<26> in1<101> in2<101> sl<52> vdd vss wl<101> / cell_PIM
XI22390 bl<58> cbl<29> in1<80> in2<80> sl<58> vdd vss wl<80> / cell_PIM
XI22389 bl<58> cbl<29> in1<81> in2<81> sl<58> vdd vss wl<81> / cell_PIM
XI21088 bl<42> cbl<21> in1<119> in2<119> sl<42> vdd vss wl<119> / cell_PIM
XI21087 bl<42> cbl<21> in1<121> in2<121> sl<42> vdd vss wl<121> / cell_PIM
XI21086 bl<42> cbl<21> in1<122> in2<122> sl<42> vdd vss wl<122> / cell_PIM
XI21085 bl<42> cbl<21> in1<120> in2<120> sl<42> vdd vss wl<120> / cell_PIM
XI21737 bl<50> cbl<25> in1<99> in2<99> sl<50> vdd vss wl<99> / cell_PIM
XI21736 bl<50> cbl<25> in1<100> in2<100> sl<50> vdd vss wl<100> / cell_PIM
XI21735 bl<50> cbl<25> in1<102> in2<102> sl<50> vdd vss wl<102> / cell_PIM
XI21734 bl<50> cbl<25> in1<103> in2<103> sl<50> vdd vss wl<103> / cell_PIM
XI22387 bl<58> cbl<29> in1<82> in2<82> sl<58> vdd vss wl<82> / cell_PIM
XI21079 bl<40> cbl<20> in1<118> in2<118> sl<40> vdd vss wl<118> / cell_PIM
XI21733 bl<50> cbl<25> in1<101> in2<101> sl<50> vdd vss wl<101> / cell_PIM
XI22382 bl<56> cbl<28> in1<80> in2<80> sl<56> vdd vss wl<80> / cell_PIM
XI22381 bl<56> cbl<28> in1<81> in2<81> sl<56> vdd vss wl<81> / cell_PIM
XI22380 bl<56> cbl<28> in1<83> in2<83> sl<56> vdd vss wl<83> / cell_PIM
XI22379 bl<56> cbl<28> in1<82> in2<82> sl<56> vdd vss wl<82> / cell_PIM
XI21727 bl<48> cbl<24> in1<100> in2<100> sl<48> vdd vss wl<100> / cell_PIM
XI21726 bl<48> cbl<24> in1<99> in2<99> sl<48> vdd vss wl<99> / cell_PIM
XI21725 bl<48> cbl<24> in1<103> in2<103> sl<48> vdd vss wl<103> / cell_PIM
XI21724 bl<48> cbl<24> in1<102> in2<102> sl<48> vdd vss wl<102> / cell_PIM
XI21078 bl<40> cbl<20> in1<119> in2<119> sl<40> vdd vss wl<119> / cell_PIM
XI21077 bl<40> cbl<20> in1<121> in2<121> sl<40> vdd vss wl<121> / cell_PIM
XI21076 bl<40> cbl<20> in1<122> in2<122> sl<40> vdd vss wl<122> / cell_PIM
XI21075 bl<40> cbl<20> in1<120> in2<120> sl<40> vdd vss wl<120> / cell_PIM
XI22374 bl<54> cbl<27> in1<80> in2<80> sl<54> vdd vss wl<80> / cell_PIM
XI21069 bl<38> cbl<19> in1<118> in2<118> sl<38> vdd vss wl<118> / cell_PIM
XI21723 bl<48> cbl<24> in1<101> in2<101> sl<48> vdd vss wl<101> / cell_PIM
XI22372 bl<54> cbl<27> in1<83> in2<83> sl<54> vdd vss wl<83> / cell_PIM
XI22371 bl<54> cbl<27> in1<82> in2<82> sl<54> vdd vss wl<82> / cell_PIM
XI21068 bl<38> cbl<19> in1<119> in2<119> sl<38> vdd vss wl<119> / cell_PIM
XI21067 bl<38> cbl<19> in1<121> in2<121> sl<38> vdd vss wl<121> / cell_PIM
XI21066 bl<38> cbl<19> in1<122> in2<122> sl<38> vdd vss wl<122> / cell_PIM
XI21065 bl<38> cbl<19> in1<120> in2<120> sl<38> vdd vss wl<120> / cell_PIM
XI21717 bl<46> cbl<23> in1<99> in2<99> sl<46> vdd vss wl<99> / cell_PIM
XI21716 bl<46> cbl<23> in1<100> in2<100> sl<46> vdd vss wl<100> / cell_PIM
XI21715 bl<46> cbl<23> in1<102> in2<102> sl<46> vdd vss wl<102> / cell_PIM
XI21714 bl<46> cbl<23> in1<103> in2<103> sl<46> vdd vss wl<103> / cell_PIM
XI22366 bl<52> cbl<26> in1<81> in2<81> sl<52> vdd vss wl<81> / cell_PIM
XI22365 bl<52> cbl<26> in1<80> in2<80> sl<52> vdd vss wl<80> / cell_PIM
XI22364 bl<52> cbl<26> in1<83> in2<83> sl<52> vdd vss wl<83> / cell_PIM
XI21059 bl<36> cbl<18> in1<119> in2<119> sl<36> vdd vss wl<119> / cell_PIM
XI21713 bl<46> cbl<23> in1<101> in2<101> sl<46> vdd vss wl<101> / cell_PIM
XI22357 bl<50> cbl<25> in1<81> in2<81> sl<50> vdd vss wl<81> / cell_PIM
XI22356 bl<50> cbl<25> in1<83> in2<83> sl<50> vdd vss wl<83> / cell_PIM
XI22355 bl<50> cbl<25> in1<82> in2<82> sl<50> vdd vss wl<82> / cell_PIM
XI21707 bl<44> cbl<22> in1<100> in2<100> sl<44> vdd vss wl<100> / cell_PIM
XI21706 bl<44> cbl<22> in1<99> in2<99> sl<44> vdd vss wl<99> / cell_PIM
XI21705 bl<44> cbl<22> in1<103> in2<103> sl<44> vdd vss wl<103> / cell_PIM
XI21704 bl<44> cbl<22> in1<102> in2<102> sl<44> vdd vss wl<102> / cell_PIM
XI21058 bl<36> cbl<18> in1<118> in2<118> sl<36> vdd vss wl<118> / cell_PIM
XI21057 bl<36> cbl<18> in1<122> in2<122> sl<36> vdd vss wl<122> / cell_PIM
XI21056 bl<36> cbl<18> in1<121> in2<121> sl<36> vdd vss wl<121> / cell_PIM
XI21055 bl<36> cbl<18> in1<120> in2<120> sl<36> vdd vss wl<120> / cell_PIM
XI21049 bl<34> cbl<17> in1<118> in2<118> sl<34> vdd vss wl<118> / cell_PIM
XI21703 bl<44> cbl<22> in1<101> in2<101> sl<44> vdd vss wl<101> / cell_PIM
XI22350 bl<48> cbl<24> in1<81> in2<81> sl<48> vdd vss wl<81> / cell_PIM
XI22349 bl<48> cbl<24> in1<80> in2<80> sl<48> vdd vss wl<80> / cell_PIM
XI21048 bl<34> cbl<17> in1<119> in2<119> sl<34> vdd vss wl<119> / cell_PIM
XI21047 bl<34> cbl<17> in1<121> in2<121> sl<34> vdd vss wl<121> / cell_PIM
XI21046 bl<34> cbl<17> in1<122> in2<122> sl<34> vdd vss wl<122> / cell_PIM
XI21045 bl<34> cbl<17> in1<120> in2<120> sl<34> vdd vss wl<120> / cell_PIM
XI21697 bl<42> cbl<21> in1<99> in2<99> sl<42> vdd vss wl<99> / cell_PIM
XI21696 bl<42> cbl<21> in1<100> in2<100> sl<42> vdd vss wl<100> / cell_PIM
XI21695 bl<42> cbl<21> in1<102> in2<102> sl<42> vdd vss wl<102> / cell_PIM
XI21694 bl<42> cbl<21> in1<103> in2<103> sl<42> vdd vss wl<103> / cell_PIM
XI22347 bl<48> cbl<24> in1<82> in2<82> sl<48> vdd vss wl<82> / cell_PIM
XI21039 bl<32> cbl<16> in1<119> in2<119> sl<32> vdd vss wl<119> / cell_PIM
XI21693 bl<42> cbl<21> in1<101> in2<101> sl<42> vdd vss wl<101> / cell_PIM
XI22342 bl<46> cbl<23> in1<80> in2<80> sl<46> vdd vss wl<80> / cell_PIM
XI22341 bl<46> cbl<23> in1<81> in2<81> sl<46> vdd vss wl<81> / cell_PIM
XI22340 bl<46> cbl<23> in1<83> in2<83> sl<46> vdd vss wl<83> / cell_PIM
XI22339 bl<46> cbl<23> in1<82> in2<82> sl<46> vdd vss wl<82> / cell_PIM
XI21687 bl<40> cbl<20> in1<99> in2<99> sl<40> vdd vss wl<99> / cell_PIM
XI21686 bl<40> cbl<20> in1<100> in2<100> sl<40> vdd vss wl<100> / cell_PIM
XI21685 bl<40> cbl<20> in1<102> in2<102> sl<40> vdd vss wl<102> / cell_PIM
XI21684 bl<40> cbl<20> in1<103> in2<103> sl<40> vdd vss wl<103> / cell_PIM
XI21038 bl<32> cbl<16> in1<118> in2<118> sl<32> vdd vss wl<118> / cell_PIM
XI21037 bl<32> cbl<16> in1<122> in2<122> sl<32> vdd vss wl<122> / cell_PIM
XI21036 bl<32> cbl<16> in1<121> in2<121> sl<32> vdd vss wl<121> / cell_PIM
XI21035 bl<32> cbl<16> in1<120> in2<120> sl<32> vdd vss wl<120> / cell_PIM
XI22334 bl<44> cbl<22> in1<81> in2<81> sl<44> vdd vss wl<81> / cell_PIM
XI21029 bl<62> cbl<31> in1<127> in2<127> sl<62> vdd vss wl<127> / cell_PIM
XI21683 bl<40> cbl<20> in1<101> in2<101> sl<40> vdd vss wl<101> / cell_PIM
XI22332 bl<44> cbl<22> in1<83> in2<83> sl<44> vdd vss wl<83> / cell_PIM
XI22331 bl<44> cbl<22> in1<82> in2<82> sl<44> vdd vss wl<82> / cell_PIM
XI21028 bl<62> cbl<31> in1<126> in2<126> sl<62> vdd vss wl<126> / cell_PIM
XI21027 bl<62> cbl<31> in1<125> in2<125> sl<62> vdd vss wl<125> / cell_PIM
XI21026 bl<62> cbl<31> in1<123> in2<123> sl<62> vdd vss wl<123> / cell_PIM
XI21025 bl<62> cbl<31> in1<124> in2<124> sl<62> vdd vss wl<124> / cell_PIM
XI21677 bl<38> cbl<19> in1<99> in2<99> sl<38> vdd vss wl<99> / cell_PIM
XI21676 bl<38> cbl<19> in1<100> in2<100> sl<38> vdd vss wl<100> / cell_PIM
XI21675 bl<38> cbl<19> in1<102> in2<102> sl<38> vdd vss wl<102> / cell_PIM
XI21674 bl<38> cbl<19> in1<103> in2<103> sl<38> vdd vss wl<103> / cell_PIM
XI22326 bl<42> cbl<21> in1<80> in2<80> sl<42> vdd vss wl<80> / cell_PIM
XI22325 bl<42> cbl<21> in1<81> in2<81> sl<42> vdd vss wl<81> / cell_PIM
XI22324 bl<42> cbl<21> in1<83> in2<83> sl<42> vdd vss wl<83> / cell_PIM
XI19282 bl<30> cbl<15> in1<103> in2<103> sl<30> vdd vss wl<103> / cell_PIM
XI19281 bl<30> cbl<15> in1<101> in2<101> sl<30> vdd vss wl<101> / cell_PIM
XI19283 bl<30> cbl<15> in1<102> in2<102> sl<30> vdd vss wl<102> / cell_PIM
XI19900 bl<16> cbl<8> in1<59> in2<59> sl<16> vdd vss wl<59> / cell_PIM
XI19899 bl<16> cbl<8> in1<58> in2<58> sl<16> vdd vss wl<58> / cell_PIM
XI20453 bl<18> cbl<9> in1<25> in2<25> sl<18> vdd vss wl<25> / cell_PIM
XI20447 bl<16> cbl<8> in1<24> in2<24> sl<16> vdd vss wl<24> / cell_PIM
XI20446 bl<16> cbl<8> in1<23> in2<23> sl<16> vdd vss wl<23> / cell_PIM
XI20445 bl<16> cbl<8> in1<22> in2<22> sl<16> vdd vss wl<22> / cell_PIM
XI20444 bl<16> cbl<8> in1<26> in2<26> sl<16> vdd vss wl<26> / cell_PIM
XI19894 bl<30> cbl<15> in1<61> in2<61> sl<30> vdd vss wl<61> / cell_PIM
XI19893 bl<30> cbl<15> in1<62> in2<62> sl<30> vdd vss wl<62> / cell_PIM
XI19275 bl<28> cbl<14> in1<100> in2<100> sl<28> vdd vss wl<100> / cell_PIM
XI19274 bl<28> cbl<14> in1<99> in2<99> sl<28> vdd vss wl<99> / cell_PIM
XI19272 bl<28> cbl<14> in1<102> in2<102> sl<28> vdd vss wl<102> / cell_PIM
XI19271 bl<28> cbl<14> in1<101> in2<101> sl<28> vdd vss wl<101> / cell_PIM
XI19273 bl<28> cbl<14> in1<103> in2<103> sl<28> vdd vss wl<103> / cell_PIM
XI19892 bl<30> cbl<15> in1<64> in2<64> sl<30> vdd vss wl<64> / cell_PIM
XI19891 bl<30> cbl<15> in1<63> in2<63> sl<30> vdd vss wl<63> / cell_PIM
XI20443 bl<16> cbl<8> in1<25> in2<25> sl<16> vdd vss wl<25> / cell_PIM
XI19265 bl<26> cbl<13> in1<99> in2<99> sl<26> vdd vss wl<99> / cell_PIM
XI19264 bl<26> cbl<13> in1<100> in2<100> sl<26> vdd vss wl<100> / cell_PIM
XI19886 bl<28> cbl<14> in1<62> in2<62> sl<28> vdd vss wl<62> / cell_PIM
XI19885 bl<28> cbl<14> in1<61> in2<61> sl<28> vdd vss wl<61> / cell_PIM
XI20437 bl<30> cbl<15> in1<27> in2<27> sl<30> vdd vss wl<27> / cell_PIM
XI20436 bl<30> cbl<15> in1<28> in2<28> sl<30> vdd vss wl<28> / cell_PIM
XI20435 bl<30> cbl<15> in1<30> in2<30> sl<30> vdd vss wl<30> / cell_PIM
XI20434 bl<30> cbl<15> in1<31> in2<31> sl<30> vdd vss wl<31> / cell_PIM
XI19262 bl<26> cbl<13> in1<103> in2<103> sl<26> vdd vss wl<103> / cell_PIM
XI19261 bl<26> cbl<13> in1<101> in2<101> sl<26> vdd vss wl<101> / cell_PIM
XI19263 bl<26> cbl<13> in1<102> in2<102> sl<26> vdd vss wl<102> / cell_PIM
XI19884 bl<28> cbl<14> in1<64> in2<64> sl<28> vdd vss wl<64> / cell_PIM
XI19883 bl<28> cbl<14> in1<63> in2<63> sl<28> vdd vss wl<63> / cell_PIM
XI20433 bl<30> cbl<15> in1<29> in2<29> sl<30> vdd vss wl<29> / cell_PIM
XI20427 bl<28> cbl<14> in1<28> in2<28> sl<28> vdd vss wl<28> / cell_PIM
XI20426 bl<28> cbl<14> in1<27> in2<27> sl<28> vdd vss wl<27> / cell_PIM
XI20425 bl<28> cbl<14> in1<31> in2<31> sl<28> vdd vss wl<31> / cell_PIM
XI20424 bl<28> cbl<14> in1<30> in2<30> sl<28> vdd vss wl<30> / cell_PIM
XI19878 bl<26> cbl<13> in1<61> in2<61> sl<26> vdd vss wl<61> / cell_PIM
XI19877 bl<26> cbl<13> in1<62> in2<62> sl<26> vdd vss wl<62> / cell_PIM
XI19255 bl<24> cbl<12> in1<99> in2<99> sl<24> vdd vss wl<99> / cell_PIM
XI19254 bl<24> cbl<12> in1<100> in2<100> sl<24> vdd vss wl<100> / cell_PIM
XI19252 bl<24> cbl<12> in1<103> in2<103> sl<24> vdd vss wl<103> / cell_PIM
XI19251 bl<24> cbl<12> in1<101> in2<101> sl<24> vdd vss wl<101> / cell_PIM
XI19253 bl<24> cbl<12> in1<102> in2<102> sl<24> vdd vss wl<102> / cell_PIM
XI19876 bl<26> cbl<13> in1<64> in2<64> sl<26> vdd vss wl<64> / cell_PIM
XI19875 bl<26> cbl<13> in1<63> in2<63> sl<26> vdd vss wl<63> / cell_PIM
XI20423 bl<28> cbl<14> in1<29> in2<29> sl<28> vdd vss wl<29> / cell_PIM
XI19245 bl<22> cbl<11> in1<99> in2<99> sl<22> vdd vss wl<99> / cell_PIM
XI19244 bl<22> cbl<11> in1<100> in2<100> sl<22> vdd vss wl<100> / cell_PIM
XI19870 bl<24> cbl<12> in1<61> in2<61> sl<24> vdd vss wl<61> / cell_PIM
XI19869 bl<24> cbl<12> in1<62> in2<62> sl<24> vdd vss wl<62> / cell_PIM
XI20417 bl<26> cbl<13> in1<27> in2<27> sl<26> vdd vss wl<27> / cell_PIM
XI20416 bl<26> cbl<13> in1<28> in2<28> sl<26> vdd vss wl<28> / cell_PIM
XI20415 bl<26> cbl<13> in1<30> in2<30> sl<26> vdd vss wl<30> / cell_PIM
XI20414 bl<26> cbl<13> in1<31> in2<31> sl<26> vdd vss wl<31> / cell_PIM
XI19242 bl<22> cbl<11> in1<103> in2<103> sl<22> vdd vss wl<103> / cell_PIM
XI19241 bl<22> cbl<11> in1<101> in2<101> sl<22> vdd vss wl<101> / cell_PIM
XI19243 bl<22> cbl<11> in1<102> in2<102> sl<22> vdd vss wl<102> / cell_PIM
XI19868 bl<24> cbl<12> in1<64> in2<64> sl<24> vdd vss wl<64> / cell_PIM
XI19867 bl<24> cbl<12> in1<63> in2<63> sl<24> vdd vss wl<63> / cell_PIM
XI20413 bl<26> cbl<13> in1<29> in2<29> sl<26> vdd vss wl<29> / cell_PIM
XI20407 bl<24> cbl<12> in1<27> in2<27> sl<24> vdd vss wl<27> / cell_PIM
XI20406 bl<24> cbl<12> in1<28> in2<28> sl<24> vdd vss wl<28> / cell_PIM
XI20405 bl<24> cbl<12> in1<30> in2<30> sl<24> vdd vss wl<30> / cell_PIM
XI20404 bl<24> cbl<12> in1<31> in2<31> sl<24> vdd vss wl<31> / cell_PIM
XI19862 bl<22> cbl<11> in1<61> in2<61> sl<22> vdd vss wl<61> / cell_PIM
XI19861 bl<22> cbl<11> in1<62> in2<62> sl<22> vdd vss wl<62> / cell_PIM
XI19235 bl<20> cbl<10> in1<100> in2<100> sl<20> vdd vss wl<100> / cell_PIM
XI19234 bl<20> cbl<10> in1<99> in2<99> sl<20> vdd vss wl<99> / cell_PIM
XI19232 bl<20> cbl<10> in1<102> in2<102> sl<20> vdd vss wl<102> / cell_PIM
XI19231 bl<20> cbl<10> in1<101> in2<101> sl<20> vdd vss wl<101> / cell_PIM
XI19233 bl<20> cbl<10> in1<103> in2<103> sl<20> vdd vss wl<103> / cell_PIM
XI19860 bl<22> cbl<11> in1<64> in2<64> sl<22> vdd vss wl<64> / cell_PIM
XI19859 bl<22> cbl<11> in1<63> in2<63> sl<22> vdd vss wl<63> / cell_PIM
XI20403 bl<24> cbl<12> in1<29> in2<29> sl<24> vdd vss wl<29> / cell_PIM
XI19225 bl<18> cbl<9> in1<99> in2<99> sl<18> vdd vss wl<99> / cell_PIM
XI19224 bl<18> cbl<9> in1<100> in2<100> sl<18> vdd vss wl<100> / cell_PIM
XI19854 bl<20> cbl<10> in1<62> in2<62> sl<20> vdd vss wl<62> / cell_PIM
XI19853 bl<20> cbl<10> in1<61> in2<61> sl<20> vdd vss wl<61> / cell_PIM
XI20397 bl<22> cbl<11> in1<27> in2<27> sl<22> vdd vss wl<27> / cell_PIM
XI20396 bl<22> cbl<11> in1<28> in2<28> sl<22> vdd vss wl<28> / cell_PIM
XI20395 bl<22> cbl<11> in1<30> in2<30> sl<22> vdd vss wl<30> / cell_PIM
XI20394 bl<22> cbl<11> in1<31> in2<31> sl<22> vdd vss wl<31> / cell_PIM
XI19222 bl<18> cbl<9> in1<103> in2<103> sl<18> vdd vss wl<103> / cell_PIM
XI19221 bl<18> cbl<9> in1<101> in2<101> sl<18> vdd vss wl<101> / cell_PIM
XI19223 bl<18> cbl<9> in1<102> in2<102> sl<18> vdd vss wl<102> / cell_PIM
XI19852 bl<20> cbl<10> in1<64> in2<64> sl<20> vdd vss wl<64> / cell_PIM
XI19851 bl<20> cbl<10> in1<63> in2<63> sl<20> vdd vss wl<63> / cell_PIM
XI20393 bl<22> cbl<11> in1<29> in2<29> sl<22> vdd vss wl<29> / cell_PIM
XI20387 bl<20> cbl<10> in1<28> in2<28> sl<20> vdd vss wl<28> / cell_PIM
XI20386 bl<20> cbl<10> in1<27> in2<27> sl<20> vdd vss wl<27> / cell_PIM
XI20385 bl<20> cbl<10> in1<31> in2<31> sl<20> vdd vss wl<31> / cell_PIM
XI20384 bl<20> cbl<10> in1<30> in2<30> sl<20> vdd vss wl<30> / cell_PIM
XI19846 bl<18> cbl<9> in1<61> in2<61> sl<18> vdd vss wl<61> / cell_PIM
XI19845 bl<18> cbl<9> in1<62> in2<62> sl<18> vdd vss wl<62> / cell_PIM
XI19215 bl<16> cbl<8> in1<100> in2<100> sl<16> vdd vss wl<100> / cell_PIM
XI19214 bl<16> cbl<8> in1<99> in2<99> sl<16> vdd vss wl<99> / cell_PIM
XI19212 bl<16> cbl<8> in1<102> in2<102> sl<16> vdd vss wl<102> / cell_PIM
XI19211 bl<16> cbl<8> in1<101> in2<101> sl<16> vdd vss wl<101> / cell_PIM
XI19213 bl<16> cbl<8> in1<103> in2<103> sl<16> vdd vss wl<103> / cell_PIM
XI19844 bl<18> cbl<9> in1<64> in2<64> sl<18> vdd vss wl<64> / cell_PIM
XI19843 bl<18> cbl<9> in1<63> in2<63> sl<18> vdd vss wl<63> / cell_PIM
XI20383 bl<20> cbl<10> in1<29> in2<29> sl<20> vdd vss wl<29> / cell_PIM
XI19206 bl<30> cbl<15> in1<104> in2<104> sl<30> vdd vss wl<104> / cell_PIM
XI19205 bl<30> cbl<15> in1<105> in2<105> sl<30> vdd vss wl<105> / cell_PIM
XI19204 bl<30> cbl<15> in1<107> in2<107> sl<30> vdd vss wl<107> / cell_PIM
XI19838 bl<16> cbl<8> in1<62> in2<62> sl<16> vdd vss wl<62> / cell_PIM
XI19837 bl<16> cbl<8> in1<61> in2<61> sl<16> vdd vss wl<61> / cell_PIM
XI20377 bl<18> cbl<9> in1<27> in2<27> sl<18> vdd vss wl<27> / cell_PIM
XI20376 bl<18> cbl<9> in1<28> in2<28> sl<18> vdd vss wl<28> / cell_PIM
XI20375 bl<18> cbl<9> in1<30> in2<30> sl<18> vdd vss wl<30> / cell_PIM
XI20374 bl<18> cbl<9> in1<31> in2<31> sl<18> vdd vss wl<31> / cell_PIM
XI17333 bl<6> cbl<3> in1<118> in2<118> sl<6> vdd vss wl<118> / cell_PIM
XI17332 bl<6> cbl<3> in1<119> in2<119> sl<6> vdd vss wl<119> / cell_PIM
XI17331 bl<6> cbl<3> in1<116> in2<116> sl<6> vdd vss wl<116> / cell_PIM
XI17983 bl<8> cbl<4> in1<105> in2<105> sl<8> vdd vss wl<105> / cell_PIM
XI17982 bl<8> cbl<4> in1<104> in2<104> sl<8> vdd vss wl<104> / cell_PIM
XI17981 bl<8> cbl<4> in1<103> in2<103> sl<8> vdd vss wl<103> / cell_PIM
XI17980 bl<8> cbl<4> in1<102> in2<102> sl<8> vdd vss wl<102> / cell_PIM
XI17979 bl<8> cbl<4> in1<101> in2<101> sl<8> vdd vss wl<101> / cell_PIM
XI18631 bl<8> cbl<4> in1<24> in2<24> sl<8> vdd vss wl<24> / cell_PIM
XI18630 bl<8> cbl<4> in1<23> in2<23> sl<8> vdd vss wl<23> / cell_PIM
XI18629 bl<8> cbl<4> in1<22> in2<22> sl<8> vdd vss wl<22> / cell_PIM
XI18628 bl<8> cbl<4> in1<21> in2<21> sl<8> vdd vss wl<21> / cell_PIM
XI18627 bl<8> cbl<4> in1<20> in2<20> sl<8> vdd vss wl<20> / cell_PIM
XI17326 bl<4> cbl<2> in1<119> in2<119> sl<4> vdd vss wl<119> / cell_PIM
XI17325 bl<4> cbl<2> in1<118> in2<118> sl<4> vdd vss wl<118> / cell_PIM
XI17324 bl<4> cbl<2> in1<117> in2<117> sl<4> vdd vss wl<117> / cell_PIM
XI17323 bl<4> cbl<2> in1<116> in2<116> sl<4> vdd vss wl<116> / cell_PIM
XI17973 bl<14> cbl<7> in1<107> in2<107> sl<14> vdd vss wl<107> / cell_PIM
XI17972 bl<14> cbl<7> in1<108> in2<108> sl<14> vdd vss wl<108> / cell_PIM
XI17971 bl<14> cbl<7> in1<109> in2<109> sl<14> vdd vss wl<109> / cell_PIM
XI17970 bl<14> cbl<7> in1<110> in2<110> sl<14> vdd vss wl<110> / cell_PIM
XI17969 bl<14> cbl<7> in1<106> in2<106> sl<14> vdd vss wl<106> / cell_PIM
XI18622 bl<14> cbl<7> in1<26> in2<26> sl<14> vdd vss wl<26> / cell_PIM
XI18621 bl<14> cbl<7> in1<27> in2<27> sl<14> vdd vss wl<27> / cell_PIM
XI18620 bl<14> cbl<7> in1<28> in2<28> sl<14> vdd vss wl<28> / cell_PIM
XI18619 bl<14> cbl<7> in1<25> in2<25> sl<14> vdd vss wl<25> / cell_PIM
XI17317 bl<6> cbl<3> in1<121> in2<121> sl<6> vdd vss wl<121> / cell_PIM
XI17316 bl<6> cbl<3> in1<122> in2<122> sl<6> vdd vss wl<122> / cell_PIM
XI17315 bl<6> cbl<3> in1<123> in2<123> sl<6> vdd vss wl<123> / cell_PIM
XI17314 bl<6> cbl<3> in1<124> in2<124> sl<6> vdd vss wl<124> / cell_PIM
XI18614 bl<12> cbl<6> in1<28> in2<28> sl<12> vdd vss wl<28> / cell_PIM
XI17313 bl<6> cbl<3> in1<120> in2<120> sl<6> vdd vss wl<120> / cell_PIM
XI17963 bl<12> cbl<6> in1<110> in2<110> sl<12> vdd vss wl<110> / cell_PIM
XI17962 bl<12> cbl<6> in1<109> in2<109> sl<12> vdd vss wl<109> / cell_PIM
XI17961 bl<12> cbl<6> in1<108> in2<108> sl<12> vdd vss wl<108> / cell_PIM
XI17960 bl<12> cbl<6> in1<107> in2<107> sl<12> vdd vss wl<107> / cell_PIM
XI17959 bl<12> cbl<6> in1<106> in2<106> sl<12> vdd vss wl<106> / cell_PIM
XI18613 bl<12> cbl<6> in1<27> in2<27> sl<12> vdd vss wl<27> / cell_PIM
XI18612 bl<12> cbl<6> in1<26> in2<26> sl<12> vdd vss wl<26> / cell_PIM
XI18611 bl<12> cbl<6> in1<25> in2<25> sl<12> vdd vss wl<25> / cell_PIM
XI18606 bl<10> cbl<5> in1<26> in2<26> sl<10> vdd vss wl<26> / cell_PIM
XI18605 bl<10> cbl<5> in1<27> in2<27> sl<10> vdd vss wl<27> / cell_PIM
XI18604 bl<10> cbl<5> in1<28> in2<28> sl<10> vdd vss wl<28> / cell_PIM
XI17307 bl<4> cbl<2> in1<124> in2<124> sl<4> vdd vss wl<124> / cell_PIM
XI17306 bl<4> cbl<2> in1<123> in2<123> sl<4> vdd vss wl<123> / cell_PIM
XI17305 bl<4> cbl<2> in1<122> in2<122> sl<4> vdd vss wl<122> / cell_PIM
XI17304 bl<4> cbl<2> in1<121> in2<121> sl<4> vdd vss wl<121> / cell_PIM
XI17303 bl<4> cbl<2> in1<120> in2<120> sl<4> vdd vss wl<120> / cell_PIM
XI17299 bl<6> cbl<3> in1<127> in2<127> sl<6> vdd vss wl<127> / cell_PIM
XI17953 bl<10> cbl<5> in1<107> in2<107> sl<10> vdd vss wl<107> / cell_PIM
XI17952 bl<10> cbl<5> in1<108> in2<108> sl<10> vdd vss wl<108> / cell_PIM
XI17951 bl<10> cbl<5> in1<109> in2<109> sl<10> vdd vss wl<109> / cell_PIM
XI17950 bl<10> cbl<5> in1<110> in2<110> sl<10> vdd vss wl<110> / cell_PIM
XI17949 bl<10> cbl<5> in1<106> in2<106> sl<10> vdd vss wl<106> / cell_PIM
XI18603 bl<10> cbl<5> in1<25> in2<25> sl<10> vdd vss wl<25> / cell_PIM
XI17298 bl<6> cbl<3> in1<126> in2<126> sl<6> vdd vss wl<126> / cell_PIM
XI17297 bl<6> cbl<3> in1<125> in2<125> sl<6> vdd vss wl<125> / cell_PIM
XI18598 bl<8> cbl<4> in1<28> in2<28> sl<8> vdd vss wl<28> / cell_PIM
XI18597 bl<8> cbl<4> in1<27> in2<27> sl<8> vdd vss wl<27> / cell_PIM
XI18596 bl<8> cbl<4> in1<26> in2<26> sl<8> vdd vss wl<26> / cell_PIM
XI18595 bl<8> cbl<4> in1<25> in2<25> sl<8> vdd vss wl<25> / cell_PIM
XI17293 bl<4> cbl<2> in1<127> in2<127> sl<4> vdd vss wl<127> / cell_PIM
XI17292 bl<4> cbl<2> in1<126> in2<126> sl<4> vdd vss wl<126> / cell_PIM
XI17291 bl<4> cbl<2> in1<125> in2<125> sl<4> vdd vss wl<125> / cell_PIM
XI17290 bl<2> cbl<1> in1<0> in2<0> sl<2> vdd vss wl<0> / cell_PIM
XI17943 bl<8> cbl<4> in1<110> in2<110> sl<8> vdd vss wl<110> / cell_PIM
XI17942 bl<8> cbl<4> in1<109> in2<109> sl<8> vdd vss wl<109> / cell_PIM
XI17941 bl<8> cbl<4> in1<108> in2<108> sl<8> vdd vss wl<108> / cell_PIM
XI17940 bl<8> cbl<4> in1<107> in2<107> sl<8> vdd vss wl<107> / cell_PIM
XI17939 bl<8> cbl<4> in1<106> in2<106> sl<8> vdd vss wl<106> / cell_PIM
XI18589 bl<14> cbl<7> in1<30> in2<30> sl<14> vdd vss wl<30> / cell_PIM
XI18588 bl<14> cbl<7> in1<31> in2<31> sl<14> vdd vss wl<31> / cell_PIM
XI18587 bl<14> cbl<7> in1<32> in2<32> sl<14> vdd vss wl<32> / cell_PIM
XI18586 bl<14> cbl<7> in1<33> in2<33> sl<14> vdd vss wl<33> / cell_PIM
XI18585 bl<14> cbl<7> in1<29> in2<29> sl<14> vdd vss wl<29> / cell_PIM
XI17288 bl<2> cbl<1> in1<4> in2<4> sl<2> vdd vss wl<4> / cell_PIM
XI17287 bl<2> cbl<1> in1<3> in2<3> sl<2> vdd vss wl<3> / cell_PIM
XI17286 bl<2> cbl<1> in1<2> in2<2> sl<2> vdd vss wl<2> / cell_PIM
XI17285 bl<2> cbl<1> in1<1> in2<1> sl<2> vdd vss wl<1> / cell_PIM
XI17933 bl<14> cbl<7> in1<112> in2<112> sl<14> vdd vss wl<112> / cell_PIM
XI17932 bl<14> cbl<7> in1<113> in2<113> sl<14> vdd vss wl<113> / cell_PIM
XI17931 bl<14> cbl<7> in1<114> in2<114> sl<14> vdd vss wl<114> / cell_PIM
XI17930 bl<14> cbl<7> in1<115> in2<115> sl<14> vdd vss wl<115> / cell_PIM
XI17929 bl<14> cbl<7> in1<111> in2<111> sl<14> vdd vss wl<111> / cell_PIM
XI18579 bl<12> cbl<6> in1<33> in2<33> sl<12> vdd vss wl<33> / cell_PIM
XI17275 bl<2> cbl<1> in1<9> in2<9> sl<2> vdd vss wl<9> / cell_PIM
XI17274 bl<2> cbl<1> in1<8> in2<8> sl<2> vdd vss wl<8> / cell_PIM
XI18578 bl<12> cbl<6> in1<32> in2<32> sl<12> vdd vss wl<32> / cell_PIM
XI18577 bl<12> cbl<6> in1<31> in2<31> sl<12> vdd vss wl<31> / cell_PIM
XI18576 bl<12> cbl<6> in1<30> in2<30> sl<12> vdd vss wl<30> / cell_PIM
XI18575 bl<12> cbl<6> in1<29> in2<29> sl<12> vdd vss wl<29> / cell_PIM
XI17273 bl<2> cbl<1> in1<7> in2<7> sl<2> vdd vss wl<7> / cell_PIM
XI17272 bl<2> cbl<1> in1<6> in2<6> sl<2> vdd vss wl<6> / cell_PIM
XI17271 bl<2> cbl<1> in1<5> in2<5> sl<2> vdd vss wl<5> / cell_PIM
XI17923 bl<12> cbl<6> in1<115> in2<115> sl<12> vdd vss wl<115> / cell_PIM
XI17922 bl<12> cbl<6> in1<114> in2<114> sl<12> vdd vss wl<114> / cell_PIM
XI17921 bl<12> cbl<6> in1<113> in2<113> sl<12> vdd vss wl<113> / cell_PIM
XI17920 bl<12> cbl<6> in1<112> in2<112> sl<12> vdd vss wl<112> / cell_PIM
XI17919 bl<12> cbl<6> in1<111> in2<111> sl<12> vdd vss wl<111> / cell_PIM
XI18569 bl<10> cbl<5> in1<30> in2<30> sl<10> vdd vss wl<30> / cell_PIM
XI18568 bl<10> cbl<5> in1<31> in2<31> sl<10> vdd vss wl<31> / cell_PIM
XI18567 bl<10> cbl<5> in1<32> in2<32> sl<10> vdd vss wl<32> / cell_PIM
XI18566 bl<10> cbl<5> in1<33> in2<33> sl<10> vdd vss wl<33> / cell_PIM
XI18565 bl<10> cbl<5> in1<29> in2<29> sl<10> vdd vss wl<29> / cell_PIM
XI17265 bl<2> cbl<1> in1<14> in2<14> sl<2> vdd vss wl<14> / cell_PIM
XI17264 bl<2> cbl<1> in1<13> in2<13> sl<2> vdd vss wl<13> / cell_PIM
XI17263 bl<2> cbl<1> in1<12> in2<12> sl<2> vdd vss wl<12> / cell_PIM
XI17262 bl<2> cbl<1> in1<11> in2<11> sl<2> vdd vss wl<11> / cell_PIM
XI17261 bl<2> cbl<1> in1<10> in2<10> sl<2> vdd vss wl<10> / cell_PIM
XI17913 bl<10> cbl<5> in1<112> in2<112> sl<10> vdd vss wl<112> / cell_PIM
XI17912 bl<10> cbl<5> in1<113> in2<113> sl<10> vdd vss wl<113> / cell_PIM
XI17911 bl<10> cbl<5> in1<114> in2<114> sl<10> vdd vss wl<114> / cell_PIM
XI17910 bl<10> cbl<5> in1<115> in2<115> sl<10> vdd vss wl<115> / cell_PIM
XI17909 bl<10> cbl<5> in1<111> in2<111> sl<10> vdd vss wl<111> / cell_PIM
XI18559 bl<8> cbl<4> in1<33> in2<33> sl<8> vdd vss wl<33> / cell_PIM
XI17255 bl<2> cbl<1> in1<19> in2<19> sl<2> vdd vss wl<19> / cell_PIM
XI17254 bl<2> cbl<1> in1<18> in2<18> sl<2> vdd vss wl<18> / cell_PIM
XI18558 bl<8> cbl<4> in1<32> in2<32> sl<8> vdd vss wl<32> / cell_PIM
XI18557 bl<8> cbl<4> in1<31> in2<31> sl<8> vdd vss wl<31> / cell_PIM
XI18556 bl<8> cbl<4> in1<30> in2<30> sl<8> vdd vss wl<30> / cell_PIM
XI18555 bl<8> cbl<4> in1<29> in2<29> sl<8> vdd vss wl<29> / cell_PIM
XI16791 bl<0> cbl<0> in1<12> in2<12> sl<0> vdd vss wl<12> / cell_PIM
XI16790 bl<0> cbl<0> in1<11> in2<11> sl<0> vdd vss wl<11> / cell_PIM
XI16788 bl<0> cbl<0> in1<9> in2<9> sl<0> vdd vss wl<9> / cell_PIM
XI16787 bl<0> cbl<0> in1<8> in2<8> sl<0> vdd vss wl<8> / cell_PIM
XI16785 bl<0> cbl<0> in1<6> in2<6> sl<0> vdd vss wl<6> / cell_PIM
XI16784 bl<0> cbl<0> in1<5> in2<5> sl<0> vdd vss wl<5> / cell_PIM
XI16782 bl<0> cbl<0> in1<3> in2<3> sl<0> vdd vss wl<3> / cell_PIM
XI16781 bl<0> cbl<0> in1<2> in2<2> sl<0> vdd vss wl<2> / cell_PIM
XI16779 bl<0> cbl<0> in1<0> in2<0> sl<0> vdd vss wl<0> / cell_PIM
XI16847 bl<0> cbl<0> in1<68> in2<68> sl<0> vdd vss wl<68> / cell_PIM
XI16845 bl<0> cbl<0> in1<66> in2<66> sl<0> vdd vss wl<66> / cell_PIM
XI16844 bl<0> cbl<0> in1<65> in2<65> sl<0> vdd vss wl<65> / cell_PIM
XI16842 bl<0> cbl<0> in1<63> in2<63> sl<0> vdd vss wl<63> / cell_PIM
XI16841 bl<0> cbl<0> in1<62> in2<62> sl<0> vdd vss wl<62> / cell_PIM
XI16839 bl<0> cbl<0> in1<60> in2<60> sl<0> vdd vss wl<60> / cell_PIM
XI16838 bl<0> cbl<0> in1<59> in2<59> sl<0> vdd vss wl<59> / cell_PIM
XI22323 bl<42> cbl<21> in1<82> in2<82> sl<42> vdd vss wl<82> / cell_PIM
XI22956 bl<48> cbl<24> in1<64> in2<64> sl<48> vdd vss wl<64> / cell_PIM
XI22955 bl<48> cbl<24> in1<63> in2<63> sl<48> vdd vss wl<63> / cell_PIM
XI23493 bl<62> cbl<31> in1<46> in2<46> sl<62> vdd vss wl<46> / cell_PIM
XI23492 bl<62> cbl<31> in1<47> in2<47> sl<62> vdd vss wl<47> / cell_PIM
XI23491 bl<62> cbl<31> in1<49> in2<49> sl<62> vdd vss wl<49> / cell_PIM
XI23490 bl<62> cbl<31> in1<50> in2<50> sl<62> vdd vss wl<50> / cell_PIM
XI23489 bl<62> cbl<31> in1<48> in2<48> sl<62> vdd vss wl<48> / cell_PIM
XI24141 bl<38> cbl<19> in1<22> in2<22> sl<38> vdd vss wl<22> / cell_PIM
XI24140 bl<38> cbl<19> in1<23> in2<23> sl<38> vdd vss wl<23> / cell_PIM
XI24139 bl<38> cbl<19> in1<24> in2<24> sl<38> vdd vss wl<24> / cell_PIM
XI24789 bl<46> cbl<23> in1<3> in2<3> sl<46> vdd vss wl<3> / cell_PIM
XI24788 bl<46> cbl<23> in1<4> in2<4> sl<46> vdd vss wl<4> / cell_PIM
XI24787 bl<46> cbl<23> in1<6> in2<6> sl<46> vdd vss wl<6> / cell_PIM
XI24786 bl<46> cbl<23> in1<7> in2<7> sl<46> vdd vss wl<7> / cell_PIM
XI24785 bl<46> cbl<23> in1<5> in2<5> sl<46> vdd vss wl<5> / cell_PIM
XI24138 bl<38> cbl<19> in1<26> in2<26> sl<38> vdd vss wl<26> / cell_PIM
XI24137 bl<38> cbl<19> in1<25> in2<25> sl<38> vdd vss wl<25> / cell_PIM
XI22950 bl<46> cbl<23> in1<61> in2<61> sl<46> vdd vss wl<61> / cell_PIM
XI22949 bl<46> cbl<23> in1<62> in2<62> sl<46> vdd vss wl<62> / cell_PIM
XI22318 bl<40> cbl<20> in1<80> in2<80> sl<40> vdd vss wl<80> / cell_PIM
XI22948 bl<46> cbl<23> in1<64> in2<64> sl<46> vdd vss wl<64> / cell_PIM
XI22947 bl<46> cbl<23> in1<63> in2<63> sl<46> vdd vss wl<63> / cell_PIM
XI23483 bl<60> cbl<30> in1<47> in2<47> sl<60> vdd vss wl<47> / cell_PIM
XI23482 bl<60> cbl<30> in1<46> in2<46> sl<60> vdd vss wl<46> / cell_PIM
XI23481 bl<60> cbl<30> in1<50> in2<50> sl<60> vdd vss wl<50> / cell_PIM
XI23480 bl<60> cbl<30> in1<49> in2<49> sl<60> vdd vss wl<49> / cell_PIM
XI23479 bl<60> cbl<30> in1<48> in2<48> sl<60> vdd vss wl<48> / cell_PIM
XI24131 bl<36> cbl<18> in1<24> in2<24> sl<36> vdd vss wl<24> / cell_PIM
XI24130 bl<36> cbl<18> in1<23> in2<23> sl<36> vdd vss wl<23> / cell_PIM
XI24129 bl<36> cbl<18> in1<22> in2<22> sl<36> vdd vss wl<22> / cell_PIM
XI24779 bl<44> cbl<22> in1<4> in2<4> sl<44> vdd vss wl<4> / cell_PIM
XI22308 bl<38> cbl<19> in1<83> in2<83> sl<38> vdd vss wl<83> / cell_PIM
XI22942 bl<44> cbl<22> in1<62> in2<62> sl<44> vdd vss wl<62> / cell_PIM
XI22941 bl<44> cbl<22> in1<61> in2<61> sl<44> vdd vss wl<61> / cell_PIM
XI24127 bl<36> cbl<18> in1<25> in2<25> sl<36> vdd vss wl<25> / cell_PIM
XI24128 bl<36> cbl<18> in1<26> in2<26> sl<36> vdd vss wl<26> / cell_PIM
XI24777 bl<44> cbl<22> in1<7> in2<7> sl<44> vdd vss wl<7> / cell_PIM
XI24776 bl<44> cbl<22> in1<6> in2<6> sl<44> vdd vss wl<6> / cell_PIM
XI24775 bl<44> cbl<22> in1<5> in2<5> sl<44> vdd vss wl<5> / cell_PIM
XI24778 bl<44> cbl<22> in1<3> in2<3> sl<44> vdd vss wl<3> / cell_PIM
XI22940 bl<44> cbl<22> in1<64> in2<64> sl<44> vdd vss wl<64> / cell_PIM
XI22939 bl<44> cbl<22> in1<63> in2<63> sl<44> vdd vss wl<63> / cell_PIM
XI23473 bl<58> cbl<29> in1<46> in2<46> sl<58> vdd vss wl<46> / cell_PIM
XI23472 bl<58> cbl<29> in1<47> in2<47> sl<58> vdd vss wl<47> / cell_PIM
XI23471 bl<58> cbl<29> in1<49> in2<49> sl<58> vdd vss wl<49> / cell_PIM
XI23470 bl<58> cbl<29> in1<50> in2<50> sl<58> vdd vss wl<50> / cell_PIM
XI23469 bl<58> cbl<29> in1<48> in2<48> sl<58> vdd vss wl<48> / cell_PIM
XI24121 bl<34> cbl<17> in1<22> in2<22> sl<34> vdd vss wl<22> / cell_PIM
XI24120 bl<34> cbl<17> in1<23> in2<23> sl<34> vdd vss wl<23> / cell_PIM
XI24119 bl<34> cbl<17> in1<24> in2<24> sl<34> vdd vss wl<24> / cell_PIM
XI24769 bl<42> cbl<21> in1<3> in2<3> sl<42> vdd vss wl<3> / cell_PIM
XI24768 bl<42> cbl<21> in1<4> in2<4> sl<42> vdd vss wl<4> / cell_PIM
XI24767 bl<42> cbl<21> in1<6> in2<6> sl<42> vdd vss wl<6> / cell_PIM
XI24766 bl<42> cbl<21> in1<7> in2<7> sl<42> vdd vss wl<7> / cell_PIM
XI24765 bl<42> cbl<21> in1<5> in2<5> sl<42> vdd vss wl<5> / cell_PIM
XI24118 bl<34> cbl<17> in1<26> in2<26> sl<34> vdd vss wl<26> / cell_PIM
XI24117 bl<34> cbl<17> in1<25> in2<25> sl<34> vdd vss wl<25> / cell_PIM
XI22934 bl<42> cbl<21> in1<61> in2<61> sl<42> vdd vss wl<61> / cell_PIM
XI22933 bl<42> cbl<21> in1<62> in2<62> sl<42> vdd vss wl<62> / cell_PIM
XI22293 bl<34> cbl<17> in1<81> in2<81> sl<34> vdd vss wl<81> / cell_PIM
XI22932 bl<42> cbl<21> in1<64> in2<64> sl<42> vdd vss wl<64> / cell_PIM
XI22931 bl<42> cbl<21> in1<63> in2<63> sl<42> vdd vss wl<63> / cell_PIM
XI23463 bl<56> cbl<28> in1<46> in2<46> sl<56> vdd vss wl<46> / cell_PIM
XI23462 bl<56> cbl<28> in1<47> in2<47> sl<56> vdd vss wl<47> / cell_PIM
XI23461 bl<56> cbl<28> in1<49> in2<49> sl<56> vdd vss wl<49> / cell_PIM
XI23460 bl<56> cbl<28> in1<50> in2<50> sl<56> vdd vss wl<50> / cell_PIM
XI23459 bl<56> cbl<28> in1<48> in2<48> sl<56> vdd vss wl<48> / cell_PIM
XI24111 bl<32> cbl<16> in1<24> in2<24> sl<32> vdd vss wl<24> / cell_PIM
XI24110 bl<32> cbl<16> in1<23> in2<23> sl<32> vdd vss wl<23> / cell_PIM
XI24109 bl<32> cbl<16> in1<22> in2<22> sl<32> vdd vss wl<22> / cell_PIM
XI24759 bl<40> cbl<20> in1<3> in2<3> sl<40> vdd vss wl<3> / cell_PIM
XI22926 bl<40> cbl<20> in1<61> in2<61> sl<40> vdd vss wl<61> / cell_PIM
XI22925 bl<40> cbl<20> in1<62> in2<62> sl<40> vdd vss wl<62> / cell_PIM
XI24107 bl<32> cbl<16> in1<25> in2<25> sl<32> vdd vss wl<25> / cell_PIM
XI24108 bl<32> cbl<16> in1<26> in2<26> sl<32> vdd vss wl<26> / cell_PIM
XI24757 bl<40> cbl<20> in1<6> in2<6> sl<40> vdd vss wl<6> / cell_PIM
XI24756 bl<40> cbl<20> in1<7> in2<7> sl<40> vdd vss wl<7> / cell_PIM
XI24755 bl<40> cbl<20> in1<5> in2<5> sl<40> vdd vss wl<5> / cell_PIM
XI24758 bl<40> cbl<20> in1<4> in2<4> sl<40> vdd vss wl<4> / cell_PIM
XI17253 bl<2> cbl<1> in1<17> in2<17> sl<2> vdd vss wl<17> / cell_PIM
XI17252 bl<2> cbl<1> in1<16> in2<16> sl<2> vdd vss wl<16> / cell_PIM
XI17251 bl<2> cbl<1> in1<15> in2<15> sl<2> vdd vss wl<15> / cell_PIM
XI17903 bl<8> cbl<4> in1<115> in2<115> sl<8> vdd vss wl<115> / cell_PIM
XI17902 bl<8> cbl<4> in1<114> in2<114> sl<8> vdd vss wl<114> / cell_PIM
XI17901 bl<8> cbl<4> in1<113> in2<113> sl<8> vdd vss wl<113> / cell_PIM
XI17900 bl<8> cbl<4> in1<112> in2<112> sl<8> vdd vss wl<112> / cell_PIM
XI17899 bl<8> cbl<4> in1<111> in2<111> sl<8> vdd vss wl<111> / cell_PIM
XI18549 bl<14> cbl<7> in1<35> in2<35> sl<14> vdd vss wl<35> / cell_PIM
XI19203 bl<30> cbl<15> in1<106> in2<106> sl<30> vdd vss wl<106> / cell_PIM
XI19836 bl<16> cbl<8> in1<64> in2<64> sl<16> vdd vss wl<64> / cell_PIM
XI19835 bl<16> cbl<8> in1<63> in2<63> sl<16> vdd vss wl<63> / cell_PIM
XI20373 bl<18> cbl<9> in1<29> in2<29> sl<18> vdd vss wl<29> / cell_PIM
XI21019 bl<60> cbl<30> in1<127> in2<127> sl<60> vdd vss wl<127> / cell_PIM
XI21673 bl<38> cbl<19> in1<101> in2<101> sl<38> vdd vss wl<101> / cell_PIM
XI22317 bl<40> cbl<20> in1<81> in2<81> sl<40> vdd vss wl<81> / cell_PIM
XI22316 bl<40> cbl<20> in1<83> in2<83> sl<40> vdd vss wl<83> / cell_PIM
XI22315 bl<40> cbl<20> in1<82> in2<82> sl<40> vdd vss wl<82> / cell_PIM
XI21667 bl<36> cbl<18> in1<100> in2<100> sl<36> vdd vss wl<100> / cell_PIM
XI21666 bl<36> cbl<18> in1<99> in2<99> sl<36> vdd vss wl<99> / cell_PIM
XI21665 bl<36> cbl<18> in1<103> in2<103> sl<36> vdd vss wl<103> / cell_PIM
XI21664 bl<36> cbl<18> in1<102> in2<102> sl<36> vdd vss wl<102> / cell_PIM
XI21018 bl<60> cbl<30> in1<126> in2<126> sl<60> vdd vss wl<126> / cell_PIM
XI21017 bl<60> cbl<30> in1<125> in2<125> sl<60> vdd vss wl<125> / cell_PIM
XI21016 bl<60> cbl<30> in1<124> in2<124> sl<60> vdd vss wl<124> / cell_PIM
XI21015 bl<60> cbl<30> in1<123> in2<123> sl<60> vdd vss wl<123> / cell_PIM
XI20367 bl<16> cbl<8> in1<28> in2<28> sl<16> vdd vss wl<28> / cell_PIM
XI20366 bl<16> cbl<8> in1<27> in2<27> sl<16> vdd vss wl<27> / cell_PIM
XI20365 bl<16> cbl<8> in1<31> in2<31> sl<16> vdd vss wl<31> / cell_PIM
XI20364 bl<16> cbl<8> in1<30> in2<30> sl<16> vdd vss wl<30> / cell_PIM
XI19829 bl<30> cbl<15> in1<65> in2<65> sl<30> vdd vss wl<65> / cell_PIM
XI19198 bl<28> cbl<14> in1<105> in2<105> sl<28> vdd vss wl<105> / cell_PIM
XI19197 bl<28> cbl<14> in1<104> in2<104> sl<28> vdd vss wl<104> / cell_PIM
XI19196 bl<28> cbl<14> in1<107> in2<107> sl<28> vdd vss wl<107> / cell_PIM
XI19195 bl<28> cbl<14> in1<106> in2<106> sl<28> vdd vss wl<106> / cell_PIM
XI18548 bl<14> cbl<7> in1<36> in2<36> sl<14> vdd vss wl<36> / cell_PIM
XI18547 bl<14> cbl<7> in1<37> in2<37> sl<14> vdd vss wl<37> / cell_PIM
XI18546 bl<14> cbl<7> in1<38> in2<38> sl<14> vdd vss wl<38> / cell_PIM
XI18545 bl<14> cbl<7> in1<34> in2<34> sl<14> vdd vss wl<34> / cell_PIM
XI17894 bl<14> cbl<7> in1<117> in2<117> sl<14> vdd vss wl<117> / cell_PIM
XI17245 bl<2> cbl<1> in1<24> in2<24> sl<2> vdd vss wl<24> / cell_PIM
XI17244 bl<2> cbl<1> in1<23> in2<23> sl<2> vdd vss wl<23> / cell_PIM
XI17243 bl<2> cbl<1> in1<22> in2<22> sl<2> vdd vss wl<22> / cell_PIM
XI17242 bl<2> cbl<1> in1<21> in2<21> sl<2> vdd vss wl<21> / cell_PIM
XI17241 bl<2> cbl<1> in1<20> in2<20> sl<2> vdd vss wl<20> / cell_PIM
XI17893 bl<14> cbl<7> in1<118> in2<118> sl<14> vdd vss wl<118> / cell_PIM
XI17892 bl<14> cbl<7> in1<119> in2<119> sl<14> vdd vss wl<119> / cell_PIM
XI17891 bl<14> cbl<7> in1<116> in2<116> sl<14> vdd vss wl<116> / cell_PIM
XI18539 bl<12> cbl<6> in1<38> in2<38> sl<12> vdd vss wl<38> / cell_PIM
XI19190 bl<26> cbl<13> in1<104> in2<104> sl<26> vdd vss wl<104> / cell_PIM
XI19189 bl<26> cbl<13> in1<105> in2<105> sl<26> vdd vss wl<105> / cell_PIM
XI19828 bl<30> cbl<15> in1<66> in2<66> sl<30> vdd vss wl<66> / cell_PIM
XI19827 bl<30> cbl<15> in1<67> in2<67> sl<30> vdd vss wl<67> / cell_PIM
XI19826 bl<30> cbl<15> in1<69> in2<69> sl<30> vdd vss wl<69> / cell_PIM
XI19825 bl<30> cbl<15> in1<68> in2<68> sl<30> vdd vss wl<68> / cell_PIM
XI20363 bl<16> cbl<8> in1<29> in2<29> sl<16> vdd vss wl<29> / cell_PIM
XI21009 bl<58> cbl<29> in1<127> in2<127> sl<58> vdd vss wl<127> / cell_PIM
XI21663 bl<36> cbl<18> in1<101> in2<101> sl<36> vdd vss wl<101> / cell_PIM
XI22310 bl<38> cbl<19> in1<80> in2<80> sl<38> vdd vss wl<80> / cell_PIM
XI22309 bl<38> cbl<19> in1<81> in2<81> sl<38> vdd vss wl<81> / cell_PIM
XI17236 bl<2> cbl<1> in1<28> in2<28> sl<2> vdd vss wl<28> / cell_PIM
XI17235 bl<2> cbl<1> in1<27> in2<27> sl<2> vdd vss wl<27> / cell_PIM
XI17234 bl<2> cbl<1> in1<26> in2<26> sl<2> vdd vss wl<26> / cell_PIM
XI17886 bl<12> cbl<6> in1<119> in2<119> sl<12> vdd vss wl<119> / cell_PIM
XI17885 bl<12> cbl<6> in1<118> in2<118> sl<12> vdd vss wl<118> / cell_PIM
XI17884 bl<12> cbl<6> in1<117> in2<117> sl<12> vdd vss wl<117> / cell_PIM
XI18538 bl<12> cbl<6> in1<37> in2<37> sl<12> vdd vss wl<37> / cell_PIM
XI18537 bl<12> cbl<6> in1<36> in2<36> sl<12> vdd vss wl<36> / cell_PIM
XI18536 bl<12> cbl<6> in1<35> in2<35> sl<12> vdd vss wl<35> / cell_PIM
XI18535 bl<12> cbl<6> in1<34> in2<34> sl<12> vdd vss wl<34> / cell_PIM
XI19187 bl<26> cbl<13> in1<106> in2<106> sl<26> vdd vss wl<106> / cell_PIM
XI19188 bl<26> cbl<13> in1<107> in2<107> sl<26> vdd vss wl<107> / cell_PIM
XI20357 bl<30> cbl<15> in1<32> in2<32> sl<30> vdd vss wl<32> / cell_PIM
XI20356 bl<30> cbl<15> in1<33> in2<33> sl<30> vdd vss wl<33> / cell_PIM
XI20355 bl<30> cbl<15> in1<35> in2<35> sl<30> vdd vss wl<35> / cell_PIM
XI20354 bl<30> cbl<15> in1<36> in2<36> sl<30> vdd vss wl<36> / cell_PIM
XI21008 bl<58> cbl<29> in1<126> in2<126> sl<58> vdd vss wl<126> / cell_PIM
XI21007 bl<58> cbl<29> in1<125> in2<125> sl<58> vdd vss wl<125> / cell_PIM
XI21006 bl<58> cbl<29> in1<123> in2<123> sl<58> vdd vss wl<123> / cell_PIM
XI21005 bl<58> cbl<29> in1<124> in2<124> sl<58> vdd vss wl<124> / cell_PIM
XI21657 bl<34> cbl<17> in1<99> in2<99> sl<34> vdd vss wl<99> / cell_PIM
XI21656 bl<34> cbl<17> in1<100> in2<100> sl<34> vdd vss wl<100> / cell_PIM
XI21655 bl<34> cbl<17> in1<102> in2<102> sl<34> vdd vss wl<102> / cell_PIM
XI21654 bl<34> cbl<17> in1<103> in2<103> sl<34> vdd vss wl<103> / cell_PIM
XI22307 bl<38> cbl<19> in1<82> in2<82> sl<38> vdd vss wl<82> / cell_PIM
XI17233 bl<2> cbl<1> in1<25> in2<25> sl<2> vdd vss wl<25> / cell_PIM
XI17883 bl<12> cbl<6> in1<116> in2<116> sl<12> vdd vss wl<116> / cell_PIM
XI18529 bl<10> cbl<5> in1<35> in2<35> sl<10> vdd vss wl<35> / cell_PIM
XI19182 bl<24> cbl<12> in1<104> in2<104> sl<24> vdd vss wl<104> / cell_PIM
XI19181 bl<24> cbl<12> in1<105> in2<105> sl<24> vdd vss wl<105> / cell_PIM
XI19180 bl<24> cbl<12> in1<107> in2<107> sl<24> vdd vss wl<107> / cell_PIM
XI19179 bl<24> cbl<12> in1<106> in2<106> sl<24> vdd vss wl<106> / cell_PIM
XI19819 bl<28> cbl<14> in1<67> in2<67> sl<28> vdd vss wl<67> / cell_PIM
XI19818 bl<28> cbl<14> in1<66> in2<66> sl<28> vdd vss wl<66> / cell_PIM
XI19817 bl<28> cbl<14> in1<65> in2<65> sl<28> vdd vss wl<65> / cell_PIM
XI20353 bl<30> cbl<15> in1<34> in2<34> sl<30> vdd vss wl<34> / cell_PIM
XI20999 bl<56> cbl<28> in1<127> in2<127> sl<56> vdd vss wl<127> / cell_PIM
XI21653 bl<34> cbl<17> in1<101> in2<101> sl<34> vdd vss wl<101> / cell_PIM
XI22302 bl<36> cbl<18> in1<81> in2<81> sl<36> vdd vss wl<81> / cell_PIM
XI22301 bl<36> cbl<18> in1<80> in2<80> sl<36> vdd vss wl<80> / cell_PIM
XI22300 bl<36> cbl<18> in1<83> in2<83> sl<36> vdd vss wl<83> / cell_PIM
XI22299 bl<36> cbl<18> in1<82> in2<82> sl<36> vdd vss wl<82> / cell_PIM
XI21647 bl<32> cbl<16> in1<100> in2<100> sl<32> vdd vss wl<100> / cell_PIM
XI21646 bl<32> cbl<16> in1<99> in2<99> sl<32> vdd vss wl<99> / cell_PIM
XI21645 bl<32> cbl<16> in1<103> in2<103> sl<32> vdd vss wl<103> / cell_PIM
XI21644 bl<32> cbl<16> in1<102> in2<102> sl<32> vdd vss wl<102> / cell_PIM
XI20998 bl<56> cbl<28> in1<126> in2<126> sl<56> vdd vss wl<126> / cell_PIM
XI20997 bl<56> cbl<28> in1<125> in2<125> sl<56> vdd vss wl<125> / cell_PIM
XI20996 bl<56> cbl<28> in1<123> in2<123> sl<56> vdd vss wl<123> / cell_PIM
XI20995 bl<56> cbl<28> in1<124> in2<124> sl<56> vdd vss wl<124> / cell_PIM
XI20347 bl<28> cbl<14> in1<33> in2<33> sl<28> vdd vss wl<33> / cell_PIM
XI20346 bl<28> cbl<14> in1<32> in2<32> sl<28> vdd vss wl<32> / cell_PIM
XI20345 bl<28> cbl<14> in1<36> in2<36> sl<28> vdd vss wl<36> / cell_PIM
XI20344 bl<28> cbl<14> in1<35> in2<35> sl<28> vdd vss wl<35> / cell_PIM
XI19816 bl<28> cbl<14> in1<69> in2<69> sl<28> vdd vss wl<69> / cell_PIM
XI19815 bl<28> cbl<14> in1<68> in2<68> sl<28> vdd vss wl<68> / cell_PIM
XI19174 bl<22> cbl<11> in1<104> in2<104> sl<22> vdd vss wl<104> / cell_PIM
XI18528 bl<10> cbl<5> in1<36> in2<36> sl<10> vdd vss wl<36> / cell_PIM
XI18527 bl<10> cbl<5> in1<37> in2<37> sl<10> vdd vss wl<37> / cell_PIM
XI18526 bl<10> cbl<5> in1<38> in2<38> sl<10> vdd vss wl<38> / cell_PIM
XI18525 bl<10> cbl<5> in1<34> in2<34> sl<10> vdd vss wl<34> / cell_PIM
XI17878 bl<10> cbl<5> in1<117> in2<117> sl<10> vdd vss wl<117> / cell_PIM
XI17877 bl<10> cbl<5> in1<118> in2<118> sl<10> vdd vss wl<118> / cell_PIM
XI17876 bl<10> cbl<5> in1<119> in2<119> sl<10> vdd vss wl<119> / cell_PIM
XI17875 bl<10> cbl<5> in1<116> in2<116> sl<10> vdd vss wl<116> / cell_PIM
XI17227 bl<2> cbl<1> in1<33> in2<33> sl<2> vdd vss wl<33> / cell_PIM
XI17226 bl<2> cbl<1> in1<32> in2<32> sl<2> vdd vss wl<32> / cell_PIM
XI17225 bl<2> cbl<1> in1<31> in2<31> sl<2> vdd vss wl<31> / cell_PIM
XI17224 bl<2> cbl<1> in1<30> in2<30> sl<2> vdd vss wl<30> / cell_PIM
XI22294 bl<34> cbl<17> in1<80> in2<80> sl<34> vdd vss wl<80> / cell_PIM
XI17223 bl<2> cbl<1> in1<29> in2<29> sl<2> vdd vss wl<29> / cell_PIM
XI17870 bl<8> cbl<4> in1<119> in2<119> sl<8> vdd vss wl<119> / cell_PIM
XI17869 bl<8> cbl<4> in1<118> in2<118> sl<8> vdd vss wl<118> / cell_PIM
XI18519 bl<8> cbl<4> in1<38> in2<38> sl<8> vdd vss wl<38> / cell_PIM
XI19172 bl<22> cbl<11> in1<107> in2<107> sl<22> vdd vss wl<107> / cell_PIM
XI19171 bl<22> cbl<11> in1<106> in2<106> sl<22> vdd vss wl<106> / cell_PIM
XI19173 bl<22> cbl<11> in1<105> in2<105> sl<22> vdd vss wl<105> / cell_PIM
XI19809 bl<26> cbl<13> in1<65> in2<65> sl<26> vdd vss wl<65> / cell_PIM
XI20343 bl<28> cbl<14> in1<34> in2<34> sl<28> vdd vss wl<34> / cell_PIM
XI20989 bl<54> cbl<27> in1<127> in2<127> sl<54> vdd vss wl<127> / cell_PIM
XI21643 bl<32> cbl<16> in1<101> in2<101> sl<32> vdd vss wl<101> / cell_PIM
XI22292 bl<34> cbl<17> in1<83> in2<83> sl<34> vdd vss wl<83> / cell_PIM
XI22291 bl<34> cbl<17> in1<82> in2<82> sl<34> vdd vss wl<82> / cell_PIM
XI17217 bl<2> cbl<1> in1<38> in2<38> sl<2> vdd vss wl<38> / cell_PIM
XI17216 bl<2> cbl<1> in1<37> in2<37> sl<2> vdd vss wl<37> / cell_PIM
XI17215 bl<2> cbl<1> in1<36> in2<36> sl<2> vdd vss wl<36> / cell_PIM
XI17214 bl<2> cbl<1> in1<35> in2<35> sl<2> vdd vss wl<35> / cell_PIM
XI17868 bl<8> cbl<4> in1<117> in2<117> sl<8> vdd vss wl<117> / cell_PIM
XI17867 bl<8> cbl<4> in1<116> in2<116> sl<8> vdd vss wl<116> / cell_PIM
XI18518 bl<8> cbl<4> in1<37> in2<37> sl<8> vdd vss wl<37> / cell_PIM
XI18517 bl<8> cbl<4> in1<36> in2<36> sl<8> vdd vss wl<36> / cell_PIM
XI18516 bl<8> cbl<4> in1<35> in2<35> sl<8> vdd vss wl<35> / cell_PIM
XI18515 bl<8> cbl<4> in1<34> in2<34> sl<8> vdd vss wl<34> / cell_PIM
XI19166 bl<20> cbl<10> in1<105> in2<105> sl<20> vdd vss wl<105> / cell_PIM
XI19165 bl<20> cbl<10> in1<104> in2<104> sl<20> vdd vss wl<104> / cell_PIM
XI19164 bl<20> cbl<10> in1<107> in2<107> sl<20> vdd vss wl<107> / cell_PIM
XI19808 bl<26> cbl<13> in1<66> in2<66> sl<26> vdd vss wl<66> / cell_PIM
XI19807 bl<26> cbl<13> in1<67> in2<67> sl<26> vdd vss wl<67> / cell_PIM
XI19806 bl<26> cbl<13> in1<69> in2<69> sl<26> vdd vss wl<69> / cell_PIM
XI19805 bl<26> cbl<13> in1<68> in2<68> sl<26> vdd vss wl<68> / cell_PIM
XI20337 bl<26> cbl<13> in1<32> in2<32> sl<26> vdd vss wl<32> / cell_PIM
XI20336 bl<26> cbl<13> in1<33> in2<33> sl<26> vdd vss wl<33> / cell_PIM
XI20335 bl<26> cbl<13> in1<35> in2<35> sl<26> vdd vss wl<35> / cell_PIM
XI20334 bl<26> cbl<13> in1<36> in2<36> sl<26> vdd vss wl<36> / cell_PIM
XI20988 bl<54> cbl<27> in1<126> in2<126> sl<54> vdd vss wl<126> / cell_PIM
XI20987 bl<54> cbl<27> in1<125> in2<125> sl<54> vdd vss wl<125> / cell_PIM
XI20986 bl<54> cbl<27> in1<123> in2<123> sl<54> vdd vss wl<123> / cell_PIM
XI20985 bl<54> cbl<27> in1<124> in2<124> sl<54> vdd vss wl<124> / cell_PIM
XI21637 bl<62> cbl<31> in1<105> in2<105> sl<62> vdd vss wl<105> / cell_PIM
XI21636 bl<62> cbl<31> in1<107> in2<107> sl<62> vdd vss wl<107> / cell_PIM
XI21635 bl<62> cbl<31> in1<106> in2<106> sl<62> vdd vss wl<106> / cell_PIM
XI21638 bl<62> cbl<31> in1<104> in2<104> sl<62> vdd vss wl<104> / cell_PIM
XI22286 bl<32> cbl<16> in1<81> in2<81> sl<32> vdd vss wl<81> / cell_PIM
XI22285 bl<32> cbl<16> in1<80> in2<80> sl<32> vdd vss wl<80> / cell_PIM
XI22284 bl<32> cbl<16> in1<83> in2<83> sl<32> vdd vss wl<83> / cell_PIM
XI16836 bl<0> cbl<0> in1<57> in2<57> sl<0> vdd vss wl<57> / cell_PIM
XI16835 bl<0> cbl<0> in1<56> in2<56> sl<0> vdd vss wl<56> / cell_PIM
XI16833 bl<0> cbl<0> in1<54> in2<54> sl<0> vdd vss wl<54> / cell_PIM
XI16832 bl<0> cbl<0> in1<53> in2<53> sl<0> vdd vss wl<53> / cell_PIM
XI16830 bl<0> cbl<0> in1<51> in2<51> sl<0> vdd vss wl<51> / cell_PIM
XI16829 bl<0> cbl<0> in1<50> in2<50> sl<0> vdd vss wl<50> / cell_PIM
XI16827 bl<0> cbl<0> in1<48> in2<48> sl<0> vdd vss wl<48> / cell_PIM
XI16826 bl<0> cbl<0> in1<47> in2<47> sl<0> vdd vss wl<47> / cell_PIM
XI22283 bl<32> cbl<16> in1<82> in2<82> sl<32> vdd vss wl<82> / cell_PIM
XI22924 bl<40> cbl<20> in1<64> in2<64> sl<40> vdd vss wl<64> / cell_PIM
XI22923 bl<40> cbl<20> in1<63> in2<63> sl<40> vdd vss wl<63> / cell_PIM
XI23453 bl<54> cbl<27> in1<46> in2<46> sl<54> vdd vss wl<46> / cell_PIM
XI23452 bl<54> cbl<27> in1<47> in2<47> sl<54> vdd vss wl<47> / cell_PIM
XI23451 bl<54> cbl<27> in1<49> in2<49> sl<54> vdd vss wl<49> / cell_PIM
XI23450 bl<54> cbl<27> in1<50> in2<50> sl<54> vdd vss wl<50> / cell_PIM
XI23449 bl<54> cbl<27> in1<48> in2<48> sl<54> vdd vss wl<48> / cell_PIM
XI24101 bl<62> cbl<31> in1<27> in2<27> sl<62> vdd vss wl<27> / cell_PIM
XI24100 bl<62> cbl<31> in1<28> in2<28> sl<62> vdd vss wl<28> / cell_PIM
XI24099 bl<62> cbl<31> in1<30> in2<30> sl<62> vdd vss wl<30> / cell_PIM
XI24749 bl<38> cbl<19> in1<3> in2<3> sl<38> vdd vss wl<3> / cell_PIM
XI24748 bl<38> cbl<19> in1<4> in2<4> sl<38> vdd vss wl<4> / cell_PIM
XI24747 bl<38> cbl<19> in1<6> in2<6> sl<38> vdd vss wl<6> / cell_PIM
XI24746 bl<38> cbl<19> in1<7> in2<7> sl<38> vdd vss wl<7> / cell_PIM
XI24745 bl<38> cbl<19> in1<5> in2<5> sl<38> vdd vss wl<5> / cell_PIM
XI24098 bl<62> cbl<31> in1<31> in2<31> sl<62> vdd vss wl<31> / cell_PIM
XI24097 bl<62> cbl<31> in1<29> in2<29> sl<62> vdd vss wl<29> / cell_PIM
XI22918 bl<38> cbl<19> in1<61> in2<61> sl<38> vdd vss wl<61> / cell_PIM
XI22917 bl<38> cbl<19> in1<62> in2<62> sl<38> vdd vss wl<62> / cell_PIM
XI22273 bl<62> cbl<31> in1<87> in2<87> sl<62> vdd vss wl<87> / cell_PIM
XI22916 bl<38> cbl<19> in1<64> in2<64> sl<38> vdd vss wl<64> / cell_PIM
XI22915 bl<38> cbl<19> in1<63> in2<63> sl<38> vdd vss wl<63> / cell_PIM
XI23443 bl<52> cbl<26> in1<47> in2<47> sl<52> vdd vss wl<47> / cell_PIM
XI23442 bl<52> cbl<26> in1<46> in2<46> sl<52> vdd vss wl<46> / cell_PIM
XI23441 bl<52> cbl<26> in1<50> in2<50> sl<52> vdd vss wl<50> / cell_PIM
XI23440 bl<52> cbl<26> in1<49> in2<49> sl<52> vdd vss wl<49> / cell_PIM
XI23439 bl<52> cbl<26> in1<48> in2<48> sl<52> vdd vss wl<48> / cell_PIM
XI24091 bl<60> cbl<30> in1<28> in2<28> sl<60> vdd vss wl<28> / cell_PIM
XI24090 bl<60> cbl<30> in1<27> in2<27> sl<60> vdd vss wl<27> / cell_PIM
XI24089 bl<60> cbl<30> in1<31> in2<31> sl<60> vdd vss wl<31> / cell_PIM
XI24739 bl<36> cbl<18> in1<4> in2<4> sl<36> vdd vss wl<4> / cell_PIM
XI22910 bl<36> cbl<18> in1<62> in2<62> sl<36> vdd vss wl<62> / cell_PIM
XI22909 bl<36> cbl<18> in1<61> in2<61> sl<36> vdd vss wl<61> / cell_PIM
XI24087 bl<60> cbl<30> in1<29> in2<29> sl<60> vdd vss wl<29> / cell_PIM
XI24088 bl<60> cbl<30> in1<30> in2<30> sl<60> vdd vss wl<30> / cell_PIM
XI24737 bl<36> cbl<18> in1<7> in2<7> sl<36> vdd vss wl<7> / cell_PIM
XI24736 bl<36> cbl<18> in1<6> in2<6> sl<36> vdd vss wl<6> / cell_PIM
XI24735 bl<36> cbl<18> in1<5> in2<5> sl<36> vdd vss wl<5> / cell_PIM
XI24738 bl<36> cbl<18> in1<3> in2<3> sl<36> vdd vss wl<3> / cell_PIM
XI17213 bl<2> cbl<1> in1<34> in2<34> sl<2> vdd vss wl<34> / cell_PIM
XI17861 bl<14> cbl<7> in1<121> in2<121> sl<14> vdd vss wl<121> / cell_PIM
XI17860 bl<14> cbl<7> in1<122> in2<122> sl<14> vdd vss wl<122> / cell_PIM
XI17859 bl<14> cbl<7> in1<123> in2<123> sl<14> vdd vss wl<123> / cell_PIM
XI18509 bl<14> cbl<7> in1<40> in2<40> sl<14> vdd vss wl<40> / cell_PIM
XI19163 bl<20> cbl<10> in1<106> in2<106> sl<20> vdd vss wl<106> / cell_PIM
XI20333 bl<26> cbl<13> in1<34> in2<34> sl<26> vdd vss wl<34> / cell_PIM
XI20979 bl<52> cbl<26> in1<127> in2<127> sl<52> vdd vss wl<127> / cell_PIM
XI21630 bl<60> cbl<30> in1<105> in2<105> sl<60> vdd vss wl<105> / cell_PIM
XI21629 bl<60> cbl<30> in1<104> in2<104> sl<60> vdd vss wl<104> / cell_PIM
XI22277 bl<62> cbl<31> in1<84> in2<84> sl<62> vdd vss wl<84> / cell_PIM
XI22276 bl<62> cbl<31> in1<85> in2<85> sl<62> vdd vss wl<85> / cell_PIM
XI22275 bl<62> cbl<31> in1<86> in2<86> sl<62> vdd vss wl<86> / cell_PIM
XI21628 bl<60> cbl<30> in1<107> in2<107> sl<60> vdd vss wl<107> / cell_PIM
XI21627 bl<60> cbl<30> in1<106> in2<106> sl<60> vdd vss wl<106> / cell_PIM
XI20978 bl<52> cbl<26> in1<126> in2<126> sl<52> vdd vss wl<126> / cell_PIM
XI20977 bl<52> cbl<26> in1<125> in2<125> sl<52> vdd vss wl<125> / cell_PIM
XI20976 bl<52> cbl<26> in1<124> in2<124> sl<52> vdd vss wl<124> / cell_PIM
XI20975 bl<52> cbl<26> in1<123> in2<123> sl<52> vdd vss wl<123> / cell_PIM
XI20327 bl<24> cbl<12> in1<32> in2<32> sl<24> vdd vss wl<32> / cell_PIM
XI20326 bl<24> cbl<12> in1<33> in2<33> sl<24> vdd vss wl<33> / cell_PIM
XI20325 bl<24> cbl<12> in1<35> in2<35> sl<24> vdd vss wl<35> / cell_PIM
XI20324 bl<24> cbl<12> in1<36> in2<36> sl<24> vdd vss wl<36> / cell_PIM
XI19799 bl<24> cbl<12> in1<65> in2<65> sl<24> vdd vss wl<65> / cell_PIM
XI19798 bl<24> cbl<12> in1<66> in2<66> sl<24> vdd vss wl<66> / cell_PIM
XI19797 bl<24> cbl<12> in1<67> in2<67> sl<24> vdd vss wl<67> / cell_PIM
XI19158 bl<18> cbl<9> in1<104> in2<104> sl<18> vdd vss wl<104> / cell_PIM
XI19157 bl<18> cbl<9> in1<105> in2<105> sl<18> vdd vss wl<105> / cell_PIM
XI19156 bl<18> cbl<9> in1<107> in2<107> sl<18> vdd vss wl<107> / cell_PIM
XI19155 bl<18> cbl<9> in1<106> in2<106> sl<18> vdd vss wl<106> / cell_PIM
XI18508 bl<14> cbl<7> in1<41> in2<41> sl<14> vdd vss wl<41> / cell_PIM
XI18507 bl<14> cbl<7> in1<42> in2<42> sl<14> vdd vss wl<42> / cell_PIM
XI18506 bl<14> cbl<7> in1<43> in2<43> sl<14> vdd vss wl<43> / cell_PIM
XI18505 bl<14> cbl<7> in1<39> in2<39> sl<14> vdd vss wl<39> / cell_PIM
XI17858 bl<14> cbl<7> in1<124> in2<124> sl<14> vdd vss wl<124> / cell_PIM
XI17857 bl<14> cbl<7> in1<120> in2<120> sl<14> vdd vss wl<120> / cell_PIM
XI17207 bl<2> cbl<1> in1<43> in2<43> sl<2> vdd vss wl<43> / cell_PIM
XI17206 bl<2> cbl<1> in1<42> in2<42> sl<2> vdd vss wl<42> / cell_PIM
XI17205 bl<2> cbl<1> in1<41> in2<41> sl<2> vdd vss wl<41> / cell_PIM
XI17204 bl<2> cbl<1> in1<40> in2<40> sl<2> vdd vss wl<40> / cell_PIM
XI22274 bl<62> cbl<31> in1<88> in2<88> sl<62> vdd vss wl<88> / cell_PIM
XI17203 bl<2> cbl<1> in1<39> in2<39> sl<2> vdd vss wl<39> / cell_PIM
XI17851 bl<12> cbl<6> in1<124> in2<124> sl<12> vdd vss wl<124> / cell_PIM
XI17850 bl<12> cbl<6> in1<123> in2<123> sl<12> vdd vss wl<123> / cell_PIM
XI17849 bl<12> cbl<6> in1<122> in2<122> sl<12> vdd vss wl<122> / cell_PIM
XI18499 bl<12> cbl<6> in1<43> in2<43> sl<12> vdd vss wl<43> / cell_PIM
XI19150 bl<16> cbl<8> in1<105> in2<105> sl<16> vdd vss wl<105> / cell_PIM
XI19149 bl<16> cbl<8> in1<104> in2<104> sl<16> vdd vss wl<104> / cell_PIM
XI19796 bl<24> cbl<12> in1<69> in2<69> sl<24> vdd vss wl<69> / cell_PIM
XI19795 bl<24> cbl<12> in1<68> in2<68> sl<24> vdd vss wl<68> / cell_PIM
XI20323 bl<24> cbl<12> in1<34> in2<34> sl<24> vdd vss wl<34> / cell_PIM
XI20969 bl<50> cbl<25> in1<127> in2<127> sl<50> vdd vss wl<127> / cell_PIM
XI21622 bl<58> cbl<29> in1<104> in2<104> sl<58> vdd vss wl<104> / cell_PIM
XI21621 bl<58> cbl<29> in1<105> in2<105> sl<58> vdd vss wl<105> / cell_PIM
XI21620 bl<58> cbl<29> in1<107> in2<107> sl<58> vdd vss wl<107> / cell_PIM
XI21619 bl<58> cbl<29> in1<106> in2<106> sl<58> vdd vss wl<106> / cell_PIM
XI17198 bl<2> cbl<1> in1<47> in2<47> sl<2> vdd vss wl<47> / cell_PIM
XI17197 bl<2> cbl<1> in1<46> in2<46> sl<2> vdd vss wl<46> / cell_PIM
XI17196 bl<2> cbl<1> in1<45> in2<45> sl<2> vdd vss wl<45> / cell_PIM
XI17195 bl<2> cbl<1> in1<44> in2<44> sl<2> vdd vss wl<44> / cell_PIM
XI17848 bl<12> cbl<6> in1<121> in2<121> sl<12> vdd vss wl<121> / cell_PIM
XI17847 bl<12> cbl<6> in1<120> in2<120> sl<12> vdd vss wl<120> / cell_PIM
XI18498 bl<12> cbl<6> in1<42> in2<42> sl<12> vdd vss wl<42> / cell_PIM
XI18497 bl<12> cbl<6> in1<41> in2<41> sl<12> vdd vss wl<41> / cell_PIM
XI18496 bl<12> cbl<6> in1<40> in2<40> sl<12> vdd vss wl<40> / cell_PIM
XI18495 bl<12> cbl<6> in1<39> in2<39> sl<12> vdd vss wl<39> / cell_PIM
XI19147 bl<16> cbl<8> in1<106> in2<106> sl<16> vdd vss wl<106> / cell_PIM
XI19148 bl<16> cbl<8> in1<107> in2<107> sl<16> vdd vss wl<107> / cell_PIM
XI19789 bl<22> cbl<11> in1<65> in2<65> sl<22> vdd vss wl<65> / cell_PIM
XI20317 bl<22> cbl<11> in1<32> in2<32> sl<22> vdd vss wl<32> / cell_PIM
XI20316 bl<22> cbl<11> in1<33> in2<33> sl<22> vdd vss wl<33> / cell_PIM
XI20315 bl<22> cbl<11> in1<35> in2<35> sl<22> vdd vss wl<35> / cell_PIM
XI20314 bl<22> cbl<11> in1<36> in2<36> sl<22> vdd vss wl<36> / cell_PIM
XI20968 bl<50> cbl<25> in1<126> in2<126> sl<50> vdd vss wl<126> / cell_PIM
XI20967 bl<50> cbl<25> in1<125> in2<125> sl<50> vdd vss wl<125> / cell_PIM
XI20966 bl<50> cbl<25> in1<123> in2<123> sl<50> vdd vss wl<123> / cell_PIM
XI20965 bl<50> cbl<25> in1<124> in2<124> sl<50> vdd vss wl<124> / cell_PIM
XI21614 bl<56> cbl<28> in1<104> in2<104> sl<56> vdd vss wl<104> / cell_PIM
XI22267 bl<60> cbl<30> in1<86> in2<86> sl<60> vdd vss wl<86> / cell_PIM
XI22266 bl<60> cbl<30> in1<85> in2<85> sl<60> vdd vss wl<85> / cell_PIM
XI22265 bl<60> cbl<30> in1<84> in2<84> sl<60> vdd vss wl<84> / cell_PIM
XI22264 bl<60> cbl<30> in1<88> in2<88> sl<60> vdd vss wl<88> / cell_PIM
XI16815 bl<0> cbl<0> in1<36> in2<36> sl<0> vdd vss wl<36> / cell_PIM
XI16824 bl<0> cbl<0> in1<45> in2<45> sl<0> vdd vss wl<45> / cell_PIM
XI22263 bl<60> cbl<30> in1<87> in2<87> sl<60> vdd vss wl<87> / cell_PIM
XI22908 bl<36> cbl<18> in1<64> in2<64> sl<36> vdd vss wl<64> / cell_PIM
XI22907 bl<36> cbl<18> in1<63> in2<63> sl<36> vdd vss wl<63> / cell_PIM
XI23433 bl<50> cbl<25> in1<46> in2<46> sl<50> vdd vss wl<46> / cell_PIM
XI23432 bl<50> cbl<25> in1<47> in2<47> sl<50> vdd vss wl<47> / cell_PIM
XI23431 bl<50> cbl<25> in1<49> in2<49> sl<50> vdd vss wl<49> / cell_PIM
XI23430 bl<50> cbl<25> in1<50> in2<50> sl<50> vdd vss wl<50> / cell_PIM
XI23429 bl<50> cbl<25> in1<48> in2<48> sl<50> vdd vss wl<48> / cell_PIM
XI24081 bl<58> cbl<29> in1<27> in2<27> sl<58> vdd vss wl<27> / cell_PIM
XI24080 bl<58> cbl<29> in1<28> in2<28> sl<58> vdd vss wl<28> / cell_PIM
XI24079 bl<58> cbl<29> in1<30> in2<30> sl<58> vdd vss wl<30> / cell_PIM
XI24729 bl<34> cbl<17> in1<3> in2<3> sl<34> vdd vss wl<3> / cell_PIM
XI22901 bl<34> cbl<17> in1<62> in2<62> sl<34> vdd vss wl<62> / cell_PIM
XI22902 bl<34> cbl<17> in1<61> in2<61> sl<34> vdd vss wl<61> / cell_PIM
XI24077 bl<58> cbl<29> in1<29> in2<29> sl<58> vdd vss wl<29> / cell_PIM
XI24078 bl<58> cbl<29> in1<31> in2<31> sl<58> vdd vss wl<31> / cell_PIM
XI24725 bl<34> cbl<17> in1<5> in2<5> sl<34> vdd vss wl<5> / cell_PIM
XI24726 bl<34> cbl<17> in1<7> in2<7> sl<34> vdd vss wl<7> / cell_PIM
XI24727 bl<34> cbl<17> in1<6> in2<6> sl<34> vdd vss wl<6> / cell_PIM
XI24728 bl<34> cbl<17> in1<4> in2<4> sl<34> vdd vss wl<4> / cell_PIM
XI17189 bl<2> cbl<1> in1<52> in2<52> sl<2> vdd vss wl<52> / cell_PIM
XI17841 bl<10> cbl<5> in1<121> in2<121> sl<10> vdd vss wl<121> / cell_PIM
XI17840 bl<10> cbl<5> in1<122> in2<122> sl<10> vdd vss wl<122> / cell_PIM
XI17839 bl<10> cbl<5> in1<123> in2<123> sl<10> vdd vss wl<123> / cell_PIM
XI18489 bl<10> cbl<5> in1<40> in2<40> sl<10> vdd vss wl<40> / cell_PIM
XI19141 bl<30> cbl<15> in1<108> in2<108> sl<30> vdd vss wl<108> / cell_PIM
XI19140 bl<30> cbl<15> in1<109> in2<109> sl<30> vdd vss wl<109> / cell_PIM
XI19139 bl<30> cbl<15> in1<110> in2<110> sl<30> vdd vss wl<110> / cell_PIM
XI19788 bl<22> cbl<11> in1<66> in2<66> sl<22> vdd vss wl<66> / cell_PIM
XI19787 bl<22> cbl<11> in1<67> in2<67> sl<22> vdd vss wl<67> / cell_PIM
XI19786 bl<22> cbl<11> in1<69> in2<69> sl<22> vdd vss wl<69> / cell_PIM
XI19785 bl<22> cbl<11> in1<68> in2<68> sl<22> vdd vss wl<68> / cell_PIM
XI20313 bl<22> cbl<11> in1<34> in2<34> sl<22> vdd vss wl<34> / cell_PIM
XI20959 bl<48> cbl<24> in1<127> in2<127> sl<48> vdd vss wl<127> / cell_PIM
XI21612 bl<56> cbl<28> in1<107> in2<107> sl<56> vdd vss wl<107> / cell_PIM
XI21611 bl<56> cbl<28> in1<106> in2<106> sl<56> vdd vss wl<106> / cell_PIM
XI21613 bl<56> cbl<28> in1<105> in2<105> sl<56> vdd vss wl<105> / cell_PIM
XI17185 bl<2> cbl<1> in1<48> in2<48> sl<2> vdd vss wl<48> / cell_PIM
XI17186 bl<2> cbl<1> in1<49> in2<49> sl<2> vdd vss wl<49> / cell_PIM
XI17187 bl<2> cbl<1> in1<50> in2<50> sl<2> vdd vss wl<50> / cell_PIM
XI17188 bl<2> cbl<1> in1<51> in2<51> sl<2> vdd vss wl<51> / cell_PIM
XI17837 bl<10> cbl<5> in1<120> in2<120> sl<10> vdd vss wl<120> / cell_PIM
XI17838 bl<10> cbl<5> in1<124> in2<124> sl<10> vdd vss wl<124> / cell_PIM
XI18485 bl<10> cbl<5> in1<39> in2<39> sl<10> vdd vss wl<39> / cell_PIM
XI18486 bl<10> cbl<5> in1<43> in2<43> sl<10> vdd vss wl<43> / cell_PIM
XI18487 bl<10> cbl<5> in1<42> in2<42> sl<10> vdd vss wl<42> / cell_PIM
XI18488 bl<10> cbl<5> in1<41> in2<41> sl<10> vdd vss wl<41> / cell_PIM
XI19137 bl<30> cbl<15> in1<111> in2<111> sl<30> vdd vss wl<111> / cell_PIM
XI19138 bl<30> cbl<15> in1<112> in2<112> sl<30> vdd vss wl<112> / cell_PIM
XI20304 bl<20> cbl<10> in1<35> in2<35> sl<20> vdd vss wl<35> / cell_PIM
XI20305 bl<20> cbl<10> in1<36> in2<36> sl<20> vdd vss wl<36> / cell_PIM
XI20306 bl<20> cbl<10> in1<32> in2<32> sl<20> vdd vss wl<32> / cell_PIM
XI20307 bl<20> cbl<10> in1<33> in2<33> sl<20> vdd vss wl<33> / cell_PIM
XI20955 bl<48> cbl<24> in1<123> in2<123> sl<48> vdd vss wl<123> / cell_PIM
XI20956 bl<48> cbl<24> in1<124> in2<124> sl<48> vdd vss wl<124> / cell_PIM
XI20957 bl<48> cbl<24> in1<125> in2<125> sl<48> vdd vss wl<125> / cell_PIM
XI20958 bl<48> cbl<24> in1<126> in2<126> sl<48> vdd vss wl<126> / cell_PIM
XI21604 bl<54> cbl<27> in1<107> in2<107> sl<54> vdd vss wl<107> / cell_PIM
XI21605 bl<54> cbl<27> in1<105> in2<105> sl<54> vdd vss wl<105> / cell_PIM
XI21606 bl<54> cbl<27> in1<104> in2<104> sl<54> vdd vss wl<104> / cell_PIM
XI22255 bl<58> cbl<29> in1<86> in2<86> sl<58> vdd vss wl<86> / cell_PIM
XI22256 bl<58> cbl<29> in1<85> in2<85> sl<58> vdd vss wl<85> / cell_PIM
XI22257 bl<58> cbl<29> in1<84> in2<84> sl<58> vdd vss wl<84> / cell_PIM
XI22254 bl<58> cbl<29> in1<88> in2<88> sl<58> vdd vss wl<88> / cell_PIM
XI16823 bl<0> cbl<0> in1<44> in2<44> sl<0> vdd vss wl<44> / cell_PIM
XI16816 bl<0> cbl<0> in1<37> in2<37> sl<0> vdd vss wl<37> / cell_PIM
XI17179 bl<2> cbl<1> in1<57> in2<57> sl<2> vdd vss wl<57> / cell_PIM
XI17831 bl<8> cbl<4> in1<124> in2<124> sl<8> vdd vss wl<124> / cell_PIM
XI17830 bl<8> cbl<4> in1<123> in2<123> sl<8> vdd vss wl<123> / cell_PIM
XI17829 bl<8> cbl<4> in1<122> in2<122> sl<8> vdd vss wl<122> / cell_PIM
XI18479 bl<8> cbl<4> in1<43> in2<43> sl<8> vdd vss wl<43> / cell_PIM
XI19131 bl<28> cbl<14> in1<110> in2<110> sl<28> vdd vss wl<110> / cell_PIM
XI19130 bl<28> cbl<14> in1<109> in2<109> sl<28> vdd vss wl<109> / cell_PIM
XI19129 bl<28> cbl<14> in1<108> in2<108> sl<28> vdd vss wl<108> / cell_PIM
XI19779 bl<20> cbl<10> in1<67> in2<67> sl<20> vdd vss wl<67> / cell_PIM
XI19778 bl<20> cbl<10> in1<66> in2<66> sl<20> vdd vss wl<66> / cell_PIM
XI19777 bl<20> cbl<10> in1<65> in2<65> sl<20> vdd vss wl<65> / cell_PIM
XI20303 bl<20> cbl<10> in1<34> in2<34> sl<20> vdd vss wl<34> / cell_PIM
XI20949 bl<46> cbl<23> in1<127> in2<127> sl<46> vdd vss wl<127> / cell_PIM
XI21603 bl<54> cbl<27> in1<106> in2<106> sl<54> vdd vss wl<106> / cell_PIM
XI22253 bl<58> cbl<29> in1<87> in2<87> sl<58> vdd vss wl<87> / cell_PIM
XI22900 bl<34> cbl<17> in1<64> in2<64> sl<34> vdd vss wl<64> / cell_PIM
XI22899 bl<34> cbl<17> in1<63> in2<63> sl<34> vdd vss wl<63> / cell_PIM
XI23423 bl<48> cbl<24> in1<47> in2<47> sl<48> vdd vss wl<47> / cell_PIM
XI23422 bl<48> cbl<24> in1<46> in2<46> sl<48> vdd vss wl<46> / cell_PIM
XI23421 bl<48> cbl<24> in1<50> in2<50> sl<48> vdd vss wl<50> / cell_PIM
XI23420 bl<48> cbl<24> in1<49> in2<49> sl<48> vdd vss wl<49> / cell_PIM
XI23419 bl<48> cbl<24> in1<48> in2<48> sl<48> vdd vss wl<48> / cell_PIM
XI24071 bl<56> cbl<28> in1<27> in2<27> sl<56> vdd vss wl<27> / cell_PIM
XI24070 bl<56> cbl<28> in1<28> in2<28> sl<56> vdd vss wl<28> / cell_PIM
XI24069 bl<56> cbl<28> in1<30> in2<30> sl<56> vdd vss wl<30> / cell_PIM
XI24719 bl<32> cbl<16> in1<4> in2<4> sl<32> vdd vss wl<4> / cell_PIM
XI16814 bl<0> cbl<0> in1<35> in2<35> sl<0> vdd vss wl<35> / cell_PIM
XI17037 bl<2> cbl<1> in1<127> in2<127> sl<2> vdd vss wl<127> / cell_PIM
XI17178 bl<2> cbl<1> in1<56> in2<56> sl<2> vdd vss wl<56> / cell_PIM
XI17177 bl<2> cbl<1> in1<55> in2<55> sl<2> vdd vss wl<55> / cell_PIM
XI17176 bl<2> cbl<1> in1<54> in2<54> sl<2> vdd vss wl<54> / cell_PIM
XI17175 bl<2> cbl<1> in1<53> in2<53> sl<2> vdd vss wl<53> / cell_PIM
XI17828 bl<8> cbl<4> in1<121> in2<121> sl<8> vdd vss wl<121> / cell_PIM
XI17827 bl<8> cbl<4> in1<120> in2<120> sl<8> vdd vss wl<120> / cell_PIM
XI18478 bl<8> cbl<4> in1<42> in2<42> sl<8> vdd vss wl<42> / cell_PIM
XI18477 bl<8> cbl<4> in1<41> in2<41> sl<8> vdd vss wl<41> / cell_PIM
XI18476 bl<8> cbl<4> in1<40> in2<40> sl<8> vdd vss wl<40> / cell_PIM
XI18475 bl<8> cbl<4> in1<39> in2<39> sl<8> vdd vss wl<39> / cell_PIM
XI19127 bl<28> cbl<14> in1<111> in2<111> sl<28> vdd vss wl<111> / cell_PIM
XI19128 bl<28> cbl<14> in1<112> in2<112> sl<28> vdd vss wl<112> / cell_PIM
XI19776 bl<20> cbl<10> in1<69> in2<69> sl<20> vdd vss wl<69> / cell_PIM
XI19775 bl<20> cbl<10> in1<68> in2<68> sl<20> vdd vss wl<68> / cell_PIM
XI20297 bl<18> cbl<9> in1<32> in2<32> sl<18> vdd vss wl<32> / cell_PIM
XI20296 bl<18> cbl<9> in1<33> in2<33> sl<18> vdd vss wl<33> / cell_PIM
XI20295 bl<18> cbl<9> in1<35> in2<35> sl<18> vdd vss wl<35> / cell_PIM
XI20294 bl<18> cbl<9> in1<36> in2<36> sl<18> vdd vss wl<36> / cell_PIM
XI20948 bl<46> cbl<23> in1<126> in2<126> sl<46> vdd vss wl<126> / cell_PIM
XI20947 bl<46> cbl<23> in1<125> in2<125> sl<46> vdd vss wl<125> / cell_PIM
XI20946 bl<46> cbl<23> in1<123> in2<123> sl<46> vdd vss wl<123> / cell_PIM
XI20945 bl<46> cbl<23> in1<124> in2<124> sl<46> vdd vss wl<124> / cell_PIM
XI21597 bl<52> cbl<26> in1<104> in2<104> sl<52> vdd vss wl<104> / cell_PIM
XI21596 bl<52> cbl<26> in1<107> in2<107> sl<52> vdd vss wl<107> / cell_PIM
XI21595 bl<52> cbl<26> in1<106> in2<106> sl<52> vdd vss wl<106> / cell_PIM
XI21598 bl<52> cbl<26> in1<105> in2<105> sl<52> vdd vss wl<105> / cell_PIM
XI22247 bl<56> cbl<28> in1<84> in2<84> sl<56> vdd vss wl<84> / cell_PIM
XI22246 bl<56> cbl<28> in1<85> in2<85> sl<56> vdd vss wl<85> / cell_PIM
XI22245 bl<56> cbl<28> in1<86> in2<86> sl<56> vdd vss wl<86> / cell_PIM
XI22244 bl<56> cbl<28> in1<88> in2<88> sl<56> vdd vss wl<88> / cell_PIM
XI22894 bl<32> cbl<16> in1<62> in2<62> sl<32> vdd vss wl<62> / cell_PIM
XI22893 bl<32> cbl<16> in1<61> in2<61> sl<32> vdd vss wl<61> / cell_PIM
XI24067 bl<56> cbl<28> in1<29> in2<29> sl<56> vdd vss wl<29> / cell_PIM
XI24068 bl<56> cbl<28> in1<31> in2<31> sl<56> vdd vss wl<31> / cell_PIM
XI24717 bl<32> cbl<16> in1<7> in2<7> sl<32> vdd vss wl<7> / cell_PIM
XI24716 bl<32> cbl<16> in1<6> in2<6> sl<32> vdd vss wl<6> / cell_PIM
XI24715 bl<32> cbl<16> in1<5> in2<5> sl<32> vdd vss wl<5> / cell_PIM
XI24718 bl<32> cbl<16> in1<3> in2<3> sl<32> vdd vss wl<3> / cell_PIM
XI16813 bl<0> cbl<0> in1<34> in2<34> sl<0> vdd vss wl<34> / cell_PIM
XI24704 bl<61> cbl<30> in1<9> in2<9> sl<61> vdd vss wl<9> / cell_PIM2
XI24054 bl<53> cbl<26> in1<31> in2<31> sl<53> vdd vss wl<31> / cell_PIM2
XI24055 bl<53> cbl<26> in1<27> in2<27> sl<53> vdd vss wl<27> / cell_PIM2
XI24056 bl<53> cbl<26> in1<28> in2<28> sl<53> vdd vss wl<28> / cell_PIM2
XI23408 bl<45> cbl<22> in1<47> in2<47> sl<45> vdd vss wl<47> / cell_PIM2
XI23405 bl<45> cbl<22> in1<49> in2<49> sl<45> vdd vss wl<49> / cell_PIM2
XI23406 bl<45> cbl<22> in1<50> in2<50> sl<45> vdd vss wl<50> / cell_PIM2
XI23407 bl<45> cbl<22> in1<46> in2<46> sl<45> vdd vss wl<46> / cell_PIM2
XI22887 bl<63> cbl<31> in1<68> in2<68> sl<63> vdd vss wl<68> / cell_PIM2
XI22888 bl<63> cbl<31> in1<67> in2<67> sl<63> vdd vss wl<67> / cell_PIM2
XI22886 bl<63> cbl<31> in1<69> in2<69> sl<63> vdd vss wl<69> / cell_PIM2
XI22238 bl<55> cbl<27> in1<88> in2<88> sl<55> vdd vss wl<88> / cell_PIM2
XI21584 bl<49> cbl<24> in1<107> in2<107> sl<49> vdd vss wl<107> / cell_PIM2
XI21585 bl<49> cbl<24> in1<104> in2<104> sl<49> vdd vss wl<104> / cell_PIM2
XI21586 bl<49> cbl<24> in1<105> in2<105> sl<49> vdd vss wl<105> / cell_PIM2
XI20934 bl<43> cbl<21> in1<127> in2<127> sl<43> vdd vss wl<127> / cell_PIM2
XI20288 bl<17> cbl<8> in1<34> in2<34> sl<17> vdd vss wl<34> / cell_PIM2
XI19764 bl<17> cbl<8> in1<67> in2<67> sl<17> vdd vss wl<67> / cell_PIM2
XI19114 bl<25> cbl<12> in1<110> in2<110> sl<25> vdd vss wl<110> / cell_PIM2
XI19115 bl<25> cbl<12> in1<109> in2<109> sl<25> vdd vss wl<109> / cell_PIM2
XI19116 bl<25> cbl<12> in1<108> in2<108> sl<25> vdd vss wl<108> / cell_PIM2
XI18464 bl<13> cbl<6> in1<45> in2<45> sl<13> vdd vss wl<45> / cell_PIM2
XI18465 bl<13> cbl<6> in1<46> in2<46> sl<13> vdd vss wl<46> / cell_PIM2
XI18466 bl<13> cbl<6> in1<47> in2<47> sl<13> vdd vss wl<47> / cell_PIM2
XI17818 bl<13> cbl<6> in1<125> in2<125> sl<13> vdd vss wl<125> / cell_PIM2
XI17814 bl<11> cbl<5> in1<127> in2<127> sl<11> vdd vss wl<127> / cell_PIM2
XI24710 bl<63> cbl<31> in1<12> in2<12> sl<63> vdd vss wl<12> / cell_PIM2
XI24711 bl<63> cbl<31> in1<11> in2<11> sl<63> vdd vss wl<11> / cell_PIM2
XI24712 bl<63> cbl<31> in1<10> in2<10> sl<63> vdd vss wl<10> / cell_PIM2
XI24713 bl<63> cbl<31> in1<9> in2<9> sl<63> vdd vss wl<9> / cell_PIM2
XI24062 bl<55> cbl<27> in1<31> in2<31> sl<55> vdd vss wl<31> / cell_PIM2
XI24063 bl<55> cbl<27> in1<30> in2<30> sl<55> vdd vss wl<30> / cell_PIM2
XI22890 bl<63> cbl<31> in1<65> in2<65> sl<63> vdd vss wl<65> / cell_PIM2
XI22889 bl<63> cbl<31> in1<66> in2<66> sl<63> vdd vss wl<66> / cell_PIM2
XI22240 bl<55> cbl<27> in1<86> in2<86> sl<55> vdd vss wl<86> / cell_PIM2
XI22241 bl<55> cbl<27> in1<85> in2<85> sl<55> vdd vss wl<85> / cell_PIM2
XI22242 bl<55> cbl<27> in1<84> in2<84> sl<55> vdd vss wl<84> / cell_PIM2
XI22239 bl<55> cbl<27> in1<87> in2<87> sl<55> vdd vss wl<87> / cell_PIM2
XI21591 bl<51> cbl<25> in1<107> in2<107> sl<51> vdd vss wl<107> / cell_PIM2
XI21592 bl<51> cbl<25> in1<106> in2<106> sl<51> vdd vss wl<106> / cell_PIM2
XI21593 bl<51> cbl<25> in1<105> in2<105> sl<51> vdd vss wl<105> / cell_PIM2
XI20940 bl<45> cbl<22> in1<123> in2<123> sl<45> vdd vss wl<123> / cell_PIM2
XI20941 bl<45> cbl<22> in1<124> in2<124> sl<45> vdd vss wl<124> / cell_PIM2
XI20942 bl<45> cbl<22> in1<125> in2<125> sl<45> vdd vss wl<125> / cell_PIM2
XI20943 bl<45> cbl<22> in1<126> in2<126> sl<45> vdd vss wl<126> / cell_PIM2
XI20290 bl<17> cbl<8> in1<36> in2<36> sl<17> vdd vss wl<36> / cell_PIM2
XI20291 bl<17> cbl<8> in1<32> in2<32> sl<17> vdd vss wl<32> / cell_PIM2
XI20292 bl<17> cbl<8> in1<33> in2<33> sl<17> vdd vss wl<33> / cell_PIM2
XI20289 bl<17> cbl<8> in1<35> in2<35> sl<17> vdd vss wl<35> / cell_PIM2
XI19770 bl<19> cbl<9> in1<69> in2<69> sl<19> vdd vss wl<69> / cell_PIM2
XI19771 bl<19> cbl<9> in1<68> in2<68> sl<19> vdd vss wl<68> / cell_PIM2
XI19772 bl<19> cbl<9> in1<67> in2<67> sl<19> vdd vss wl<67> / cell_PIM2
XI19122 bl<27> cbl<13> in1<112> in2<112> sl<27> vdd vss wl<112> / cell_PIM2
XI19123 bl<27> cbl<13> in1<111> in2<111> sl<27> vdd vss wl<111> / cell_PIM2
XI18471 bl<15> cbl<7> in1<47> in2<47> sl<15> vdd vss wl<47> / cell_PIM2
XI18472 bl<15> cbl<7> in1<46> in2<46> sl<15> vdd vss wl<46> / cell_PIM2
XI18473 bl<15> cbl<7> in1<45> in2<45> sl<15> vdd vss wl<45> / cell_PIM2
XI17820 bl<13> cbl<6> in1<127> in2<127> sl<13> vdd vss wl<127> / cell_PIM2
XI17819 bl<13> cbl<6> in1<126> in2<126> sl<13> vdd vss wl<126> / cell_PIM2
XI17170 bl<3> cbl<1> in1<58> in2<58> sl<3> vdd vss wl<58> / cell_PIM2
XI17171 bl<3> cbl<1> in1<59> in2<59> sl<3> vdd vss wl<59> / cell_PIM2
XI17172 bl<3> cbl<1> in1<60> in2<60> sl<3> vdd vss wl<60> / cell_PIM2
XI17173 bl<3> cbl<1> in1<61> in2<61> sl<3> vdd vss wl<61> / cell_PIM2
XI17162 bl<3> cbl<1> in1<65> in2<65> sl<3> vdd vss wl<65> / cell_PIM2
XI17153 bl<3> cbl<1> in1<70> in2<70> sl<3> vdd vss wl<70> / cell_PIM2
XI17144 bl<3> cbl<1> in1<74> in2<74> sl<3> vdd vss wl<74> / cell_PIM2
XI17135 bl<3> cbl<1> in1<80> in2<80> sl<3> vdd vss wl<80> / cell_PIM2
XI17132 bl<3> cbl<1> in1<77> in2<77> sl<3> vdd vss wl<77> / cell_PIM2
XI17126 bl<3> cbl<1> in1<86> in2<86> sl<3> vdd vss wl<86> / cell_PIM2
XI17123 bl<3> cbl<1> in1<83> in2<83> sl<3> vdd vss wl<83> / cell_PIM2
XI17114 bl<3> cbl<1> in1<89> in2<89> sl<3> vdd vss wl<89> / cell_PIM2
XI17105 bl<3> cbl<1> in1<94> in2<94> sl<3> vdd vss wl<94> / cell_PIM2
XI17096 bl<3> cbl<1> in1<98> in2<98> sl<3> vdd vss wl<98> / cell_PIM2
XI17087 bl<3> cbl<1> in1<104> in2<104> sl<3> vdd vss wl<104> / cell_PIM2
XI17084 bl<3> cbl<1> in1<101> in2<101> sl<3> vdd vss wl<101> / cell_PIM2
XI17078 bl<3> cbl<1> in1<110> in2<110> sl<3> vdd vss wl<110> / cell_PIM2
XI17075 bl<3> cbl<1> in1<107> in2<107> sl<3> vdd vss wl<107> / cell_PIM2
XI17066 bl<3> cbl<1> in1<113> in2<113> sl<3> vdd vss wl<113> / cell_PIM2
XI17057 bl<3> cbl<1> in1<118> in2<118> sl<3> vdd vss wl<118> / cell_PIM2
XI17048 bl<3> cbl<1> in1<122> in2<122> sl<3> vdd vss wl<122> / cell_PIM2
XI17039 bl<3> cbl<1> in1<126> in2<126> sl<3> vdd vss wl<126> / cell_PIM2
XI17032 bl<1> cbl<0> in1<125> in2<125> sl<1> vdd vss wl<125> / cell_PIM2
XI17029 bl<1> cbl<0> in1<122> in2<122> sl<1> vdd vss wl<122> / cell_PIM2
XI17026 bl<1> cbl<0> in1<119> in2<119> sl<1> vdd vss wl<119> / cell_PIM2
XI17023 bl<1> cbl<0> in1<116> in2<116> sl<1> vdd vss wl<116> / cell_PIM2
XI17020 bl<1> cbl<0> in1<113> in2<113> sl<1> vdd vss wl<113> / cell_PIM2
XI17017 bl<1> cbl<0> in1<110> in2<110> sl<1> vdd vss wl<110> / cell_PIM2
XI17014 bl<1> cbl<0> in1<107> in2<107> sl<1> vdd vss wl<107> / cell_PIM2
XI17011 bl<1> cbl<0> in1<104> in2<104> sl<1> vdd vss wl<104> / cell_PIM2
XI17008 bl<1> cbl<0> in1<101> in2<101> sl<1> vdd vss wl<101> / cell_PIM2
XI17005 bl<1> cbl<0> in1<98> in2<98> sl<1> vdd vss wl<98> / cell_PIM2
XI17002 bl<1> cbl<0> in1<95> in2<95> sl<1> vdd vss wl<95> / cell_PIM2
XI16999 bl<1> cbl<0> in1<92> in2<92> sl<1> vdd vss wl<92> / cell_PIM2
XI16996 bl<1> cbl<0> in1<89> in2<89> sl<1> vdd vss wl<89> / cell_PIM2
XI16993 bl<1> cbl<0> in1<86> in2<86> sl<1> vdd vss wl<86> / cell_PIM2
XI16990 bl<1> cbl<0> in1<83> in2<83> sl<1> vdd vss wl<83> / cell_PIM2
XI16987 bl<1> cbl<0> in1<80> in2<80> sl<1> vdd vss wl<80> / cell_PIM2
XI16984 bl<1> cbl<0> in1<77> in2<77> sl<1> vdd vss wl<77> / cell_PIM2
XI16981 bl<1> cbl<0> in1<74> in2<74> sl<1> vdd vss wl<74> / cell_PIM2
XI16978 bl<1> cbl<0> in1<71> in2<71> sl<1> vdd vss wl<71> / cell_PIM2
XI16975 bl<1> cbl<0> in1<68> in2<68> sl<1> vdd vss wl<68> / cell_PIM2
XI16972 bl<1> cbl<0> in1<65> in2<65> sl<1> vdd vss wl<65> / cell_PIM2
XI16969 bl<1> cbl<0> in1<62> in2<62> sl<1> vdd vss wl<62> / cell_PIM2
XI16966 bl<1> cbl<0> in1<59> in2<59> sl<1> vdd vss wl<59> / cell_PIM2
XI16963 bl<1> cbl<0> in1<56> in2<56> sl<1> vdd vss wl<56> / cell_PIM2
XI16960 bl<1> cbl<0> in1<53> in2<53> sl<1> vdd vss wl<53> / cell_PIM2
XI16957 bl<1> cbl<0> in1<50> in2<50> sl<1> vdd vss wl<50> / cell_PIM2
XI16954 bl<1> cbl<0> in1<47> in2<47> sl<1> vdd vss wl<47> / cell_PIM2
XI16951 bl<1> cbl<0> in1<44> in2<44> sl<1> vdd vss wl<44> / cell_PIM2
XI16948 bl<1> cbl<0> in1<41> in2<41> sl<1> vdd vss wl<41> / cell_PIM2
XI16945 bl<1> cbl<0> in1<38> in2<38> sl<1> vdd vss wl<38> / cell_PIM2
XI16942 bl<1> cbl<0> in1<35> in2<35> sl<1> vdd vss wl<35> / cell_PIM2
XI16939 bl<1> cbl<0> in1<32> in2<32> sl<1> vdd vss wl<32> / cell_PIM2
XI16936 bl<1> cbl<0> in1<29> in2<29> sl<1> vdd vss wl<29> / cell_PIM2
XI16933 bl<1> cbl<0> in1<26> in2<26> sl<1> vdd vss wl<26> / cell_PIM2
XI16930 bl<1> cbl<0> in1<23> in2<23> sl<1> vdd vss wl<23> / cell_PIM2
XI16927 bl<1> cbl<0> in1<20> in2<20> sl<1> vdd vss wl<20> / cell_PIM2
XI16924 bl<1> cbl<0> in1<17> in2<17> sl<1> vdd vss wl<17> / cell_PIM2
XI16921 bl<1> cbl<0> in1<14> in2<14> sl<1> vdd vss wl<14> / cell_PIM2
XI16918 bl<1> cbl<0> in1<11> in2<11> sl<1> vdd vss wl<11> / cell_PIM2
XI16915 bl<1> cbl<0> in1<8> in2<8> sl<1> vdd vss wl<8> / cell_PIM2
XI16912 bl<1> cbl<0> in1<5> in2<5> sl<1> vdd vss wl<5> / cell_PIM2
XI16909 bl<1> cbl<0> in1<2> in2<2> sl<1> vdd vss wl<2> / cell_PIM2
XI17164 bl<3> cbl<1> in1<67> in2<67> sl<3> vdd vss wl<67> / cell_PIM2
XI17163 bl<3> cbl<1> in1<66> in2<66> sl<3> vdd vss wl<66> / cell_PIM2
XI17161 bl<3> cbl<1> in1<64> in2<64> sl<3> vdd vss wl<64> / cell_PIM2
XI17160 bl<3> cbl<1> in1<63> in2<63> sl<3> vdd vss wl<63> / cell_PIM2
XI17154 bl<3> cbl<1> in1<71> in2<71> sl<3> vdd vss wl<71> / cell_PIM2
XI17152 bl<3> cbl<1> in1<69> in2<69> sl<3> vdd vss wl<69> / cell_PIM2
XI17151 bl<3> cbl<1> in1<68> in2<68> sl<3> vdd vss wl<68> / cell_PIM2
XI17146 bl<3> cbl<1> in1<76> in2<76> sl<3> vdd vss wl<76> / cell_PIM2
XI17145 bl<3> cbl<1> in1<75> in2<75> sl<3> vdd vss wl<75> / cell_PIM2
XI17143 bl<3> cbl<1> in1<73> in2<73> sl<3> vdd vss wl<73> / cell_PIM2
XI17142 bl<3> cbl<1> in1<72> in2<72> sl<3> vdd vss wl<72> / cell_PIM2
XI17136 bl<3> cbl<1> in1<81> in2<81> sl<3> vdd vss wl<81> / cell_PIM2
XI17134 bl<3> cbl<1> in1<79> in2<79> sl<3> vdd vss wl<79> / cell_PIM2
XI17133 bl<3> cbl<1> in1<78> in2<78> sl<3> vdd vss wl<78> / cell_PIM2
XI17125 bl<3> cbl<1> in1<85> in2<85> sl<3> vdd vss wl<85> / cell_PIM2
XI17124 bl<3> cbl<1> in1<84> in2<84> sl<3> vdd vss wl<84> / cell_PIM2
XI17122 bl<3> cbl<1> in1<82> in2<82> sl<3> vdd vss wl<82> / cell_PIM2
XI17116 bl<3> cbl<1> in1<91> in2<91> sl<3> vdd vss wl<91> / cell_PIM2
XI17115 bl<3> cbl<1> in1<90> in2<90> sl<3> vdd vss wl<90> / cell_PIM2
XI17113 bl<3> cbl<1> in1<88> in2<88> sl<3> vdd vss wl<88> / cell_PIM2
XI17112 bl<3> cbl<1> in1<87> in2<87> sl<3> vdd vss wl<87> / cell_PIM2
XI17106 bl<3> cbl<1> in1<95> in2<95> sl<3> vdd vss wl<95> / cell_PIM2
XI17104 bl<3> cbl<1> in1<93> in2<93> sl<3> vdd vss wl<93> / cell_PIM2
XI17103 bl<3> cbl<1> in1<92> in2<92> sl<3> vdd vss wl<92> / cell_PIM2
XI17098 bl<3> cbl<1> in1<100> in2<100> sl<3> vdd vss wl<100> / cell_PIM2
XI17097 bl<3> cbl<1> in1<99> in2<99> sl<3> vdd vss wl<99> / cell_PIM2
XI17095 bl<3> cbl<1> in1<97> in2<97> sl<3> vdd vss wl<97> / cell_PIM2
XI17094 bl<3> cbl<1> in1<96> in2<96> sl<3> vdd vss wl<96> / cell_PIM2
XI17088 bl<3> cbl<1> in1<105> in2<105> sl<3> vdd vss wl<105> / cell_PIM2
XI17086 bl<3> cbl<1> in1<103> in2<103> sl<3> vdd vss wl<103> / cell_PIM2
XI17085 bl<3> cbl<1> in1<102> in2<102> sl<3> vdd vss wl<102> / cell_PIM2
XI17077 bl<3> cbl<1> in1<109> in2<109> sl<3> vdd vss wl<109> / cell_PIM2
XI17076 bl<3> cbl<1> in1<108> in2<108> sl<3> vdd vss wl<108> / cell_PIM2
XI17074 bl<3> cbl<1> in1<106> in2<106> sl<3> vdd vss wl<106> / cell_PIM2
XI17068 bl<3> cbl<1> in1<115> in2<115> sl<3> vdd vss wl<115> / cell_PIM2
XI17067 bl<3> cbl<1> in1<114> in2<114> sl<3> vdd vss wl<114> / cell_PIM2
XI17065 bl<3> cbl<1> in1<112> in2<112> sl<3> vdd vss wl<112> / cell_PIM2
XI17064 bl<3> cbl<1> in1<111> in2<111> sl<3> vdd vss wl<111> / cell_PIM2
XI17058 bl<3> cbl<1> in1<119> in2<119> sl<3> vdd vss wl<119> / cell_PIM2
XI17056 bl<3> cbl<1> in1<117> in2<117> sl<3> vdd vss wl<117> / cell_PIM2
XI17055 bl<3> cbl<1> in1<116> in2<116> sl<3> vdd vss wl<116> / cell_PIM2
XI17050 bl<3> cbl<1> in1<124> in2<124> sl<3> vdd vss wl<124> / cell_PIM2
XI17049 bl<3> cbl<1> in1<123> in2<123> sl<3> vdd vss wl<123> / cell_PIM2
XI17047 bl<3> cbl<1> in1<121> in2<121> sl<3> vdd vss wl<121> / cell_PIM2
XI17046 bl<3> cbl<1> in1<120> in2<120> sl<3> vdd vss wl<120> / cell_PIM2
XI17040 bl<3> cbl<1> in1<127> in2<127> sl<3> vdd vss wl<127> / cell_PIM2
XI17038 bl<3> cbl<1> in1<125> in2<125> sl<3> vdd vss wl<125> / cell_PIM2
XI17034 bl<1> cbl<0> in1<127> in2<127> sl<1> vdd vss wl<127> / cell_PIM2
XI17033 bl<1> cbl<0> in1<126> in2<126> sl<1> vdd vss wl<126> / cell_PIM2
XI17031 bl<1> cbl<0> in1<124> in2<124> sl<1> vdd vss wl<124> / cell_PIM2
XI17030 bl<1> cbl<0> in1<123> in2<123> sl<1> vdd vss wl<123> / cell_PIM2
XI17028 bl<1> cbl<0> in1<121> in2<121> sl<1> vdd vss wl<121> / cell_PIM2
XI17027 bl<1> cbl<0> in1<120> in2<120> sl<1> vdd vss wl<120> / cell_PIM2
XI17025 bl<1> cbl<0> in1<118> in2<118> sl<1> vdd vss wl<118> / cell_PIM2
XI17024 bl<1> cbl<0> in1<117> in2<117> sl<1> vdd vss wl<117> / cell_PIM2
XI17022 bl<1> cbl<0> in1<115> in2<115> sl<1> vdd vss wl<115> / cell_PIM2
XI17021 bl<1> cbl<0> in1<114> in2<114> sl<1> vdd vss wl<114> / cell_PIM2
XI17019 bl<1> cbl<0> in1<112> in2<112> sl<1> vdd vss wl<112> / cell_PIM2
XI17018 bl<1> cbl<0> in1<111> in2<111> sl<1> vdd vss wl<111> / cell_PIM2
XI17016 bl<1> cbl<0> in1<109> in2<109> sl<1> vdd vss wl<109> / cell_PIM2
XI17015 bl<1> cbl<0> in1<108> in2<108> sl<1> vdd vss wl<108> / cell_PIM2
XI17013 bl<1> cbl<0> in1<106> in2<106> sl<1> vdd vss wl<106> / cell_PIM2
XI17012 bl<1> cbl<0> in1<105> in2<105> sl<1> vdd vss wl<105> / cell_PIM2
XI17010 bl<1> cbl<0> in1<103> in2<103> sl<1> vdd vss wl<103> / cell_PIM2
XI17009 bl<1> cbl<0> in1<102> in2<102> sl<1> vdd vss wl<102> / cell_PIM2
XI17007 bl<1> cbl<0> in1<100> in2<100> sl<1> vdd vss wl<100> / cell_PIM2
XI17006 bl<1> cbl<0> in1<99> in2<99> sl<1> vdd vss wl<99> / cell_PIM2
XI17004 bl<1> cbl<0> in1<97> in2<97> sl<1> vdd vss wl<97> / cell_PIM2
XI17003 bl<1> cbl<0> in1<96> in2<96> sl<1> vdd vss wl<96> / cell_PIM2
XI17001 bl<1> cbl<0> in1<94> in2<94> sl<1> vdd vss wl<94> / cell_PIM2
XI17000 bl<1> cbl<0> in1<93> in2<93> sl<1> vdd vss wl<93> / cell_PIM2
XI16998 bl<1> cbl<0> in1<91> in2<91> sl<1> vdd vss wl<91> / cell_PIM2
XI16997 bl<1> cbl<0> in1<90> in2<90> sl<1> vdd vss wl<90> / cell_PIM2
XI16995 bl<1> cbl<0> in1<88> in2<88> sl<1> vdd vss wl<88> / cell_PIM2
XI16994 bl<1> cbl<0> in1<87> in2<87> sl<1> vdd vss wl<87> / cell_PIM2
XI16992 bl<1> cbl<0> in1<85> in2<85> sl<1> vdd vss wl<85> / cell_PIM2
XI16991 bl<1> cbl<0> in1<84> in2<84> sl<1> vdd vss wl<84> / cell_PIM2
XI16989 bl<1> cbl<0> in1<82> in2<82> sl<1> vdd vss wl<82> / cell_PIM2
XI16988 bl<1> cbl<0> in1<81> in2<81> sl<1> vdd vss wl<81> / cell_PIM2
XI16986 bl<1> cbl<0> in1<79> in2<79> sl<1> vdd vss wl<79> / cell_PIM2
XI16985 bl<1> cbl<0> in1<78> in2<78> sl<1> vdd vss wl<78> / cell_PIM2
XI16983 bl<1> cbl<0> in1<76> in2<76> sl<1> vdd vss wl<76> / cell_PIM2
XI16982 bl<1> cbl<0> in1<75> in2<75> sl<1> vdd vss wl<75> / cell_PIM2
XI16980 bl<1> cbl<0> in1<73> in2<73> sl<1> vdd vss wl<73> / cell_PIM2
XI16979 bl<1> cbl<0> in1<72> in2<72> sl<1> vdd vss wl<72> / cell_PIM2
XI16977 bl<1> cbl<0> in1<70> in2<70> sl<1> vdd vss wl<70> / cell_PIM2
XI16976 bl<1> cbl<0> in1<69> in2<69> sl<1> vdd vss wl<69> / cell_PIM2
XI16974 bl<1> cbl<0> in1<67> in2<67> sl<1> vdd vss wl<67> / cell_PIM2
XI16973 bl<1> cbl<0> in1<66> in2<66> sl<1> vdd vss wl<66> / cell_PIM2
XI24703 bl<61> cbl<30> in1<8> in2<8> sl<61> vdd vss wl<8> / cell_PIM2
XI24693 bl<59> cbl<29> in1<9> in2<9> sl<59> vdd vss wl<9> / cell_PIM2
XI24683 bl<57> cbl<28> in1<9> in2<9> sl<57> vdd vss wl<9> / cell_PIM2
XI24673 bl<55> cbl<27> in1<9> in2<9> sl<55> vdd vss wl<9> / cell_PIM2
XI24663 bl<53> cbl<26> in1<8> in2<8> sl<53> vdd vss wl<8> / cell_PIM2
XI24653 bl<51> cbl<25> in1<9> in2<9> sl<51> vdd vss wl<9> / cell_PIM2
XI24643 bl<49> cbl<24> in1<8> in2<8> sl<49> vdd vss wl<8> / cell_PIM2
XI24633 bl<47> cbl<23> in1<9> in2<9> sl<47> vdd vss wl<9> / cell_PIM2
XI24623 bl<45> cbl<22> in1<8> in2<8> sl<45> vdd vss wl<8> / cell_PIM2
XI24613 bl<43> cbl<21> in1<9> in2<9> sl<43> vdd vss wl<9> / cell_PIM2
XI24603 bl<41> cbl<20> in1<9> in2<9> sl<41> vdd vss wl<9> / cell_PIM2
XI24593 bl<39> cbl<19> in1<9> in2<9> sl<39> vdd vss wl<9> / cell_PIM2
XI24583 bl<37> cbl<18> in1<8> in2<8> sl<37> vdd vss wl<8> / cell_PIM2
XI25228 vss vss vdd vdd vss vdd vss vss / cell_PIM2
XI25227 vss vss in1<0> in2<0> vss vdd vss wl<0> / cell_PIM2
XI25226 vss vss in1<1> in2<1> vss vdd vss wl<1> / cell_PIM2
XI25225 vss vss in1<2> in2<2> vss vdd vss wl<2> / cell_PIM2
XI25224 vss vss in1<4> in2<4> vss vdd vss wl<4> / cell_PIM2
XI24573 bl<35> cbl<17> in1<9> in2<9> sl<35> vdd vss wl<9> / cell_PIM2
XI25222 vss vss in1<5> in2<5> vss vdd vss wl<5> / cell_PIM2
XI25221 vss vss in1<6> in2<6> vss vdd vss wl<6> / cell_PIM2
XI25220 vss vss in1<7> in2<7> vss vdd vss wl<7> / cell_PIM2
XI25219 vss vss in1<8> in2<8> vss vdd vss wl<8> / cell_PIM2
XI25223 vss vss in1<3> in2<3> vss vdd vss wl<3> / cell_PIM2
XI25217 vss vss in1<10> in2<10> vss vdd vss wl<10> / cell_PIM2
XI25216 vss vss in1<11> in2<11> vss vdd vss wl<11> / cell_PIM2
XI25215 vss vss in1<12> in2<12> vss vdd vss wl<12> / cell_PIM2
XI25214 vss vss in1<13> in2<13> vss vdd vss wl<13> / cell_PIM2
XI25218 vss vss in1<9> in2<9> vss vdd vss wl<9> / cell_PIM2
XI24563 bl<33> cbl<16> in1<8> in2<8> sl<33> vdd vss wl<8> / cell_PIM2
XI25212 vss vss in1<15> in2<15> vss vdd vss wl<15> / cell_PIM2
XI25211 vss vss in1<16> in2<16> vss vdd vss wl<16> / cell_PIM2
XI25210 vss vss in1<17> in2<17> vss vdd vss wl<17> / cell_PIM2
XI25209 vss vss in1<18> in2<18> vss vdd vss wl<18> / cell_PIM2
XI25213 vss vss in1<14> in2<14> vss vdd vss wl<14> / cell_PIM2
XI25208 vss vss in1<19> in2<19> vss vdd vss wl<19> / cell_PIM2
XI25207 vss vss in1<20> in2<20> vss vdd vss wl<20> / cell_PIM2
XI25206 vss vss in1<21> in2<21> vss vdd vss wl<21> / cell_PIM2
XI25205 vss vss in1<22> in2<22> vss vdd vss wl<22> / cell_PIM2
XI25204 vss vss in1<23> in2<23> vss vdd vss wl<23> / cell_PIM2
XI24553 bl<63> cbl<31> in1<14> in2<14> sl<63> vdd vss wl<14> / cell_PIM2
XI25202 vss vss in1<25> in2<25> vss vdd vss wl<25> / cell_PIM2
XI25201 vss vss in1<26> in2<26> vss vdd vss wl<26> / cell_PIM2
XI25200 vss vss in1<27> in2<27> vss vdd vss wl<27> / cell_PIM2
XI25199 vss vss in1<28> in2<28> vss vdd vss wl<28> / cell_PIM2
XI25203 vss vss in1<24> in2<24> vss vdd vss wl<24> / cell_PIM2
XI25197 vss vss in1<30> in2<30> vss vdd vss wl<30> / cell_PIM2
XI25196 vss vss in1<31> in2<31> vss vdd vss wl<31> / cell_PIM2
XI25195 vss vss in1<32> in2<32> vss vdd vss wl<32> / cell_PIM2
XI25194 vss vss in1<33> in2<33> vss vdd vss wl<33> / cell_PIM2
XI25198 vss vss in1<29> in2<29> vss vdd vss wl<29> / cell_PIM2
XI24543 bl<61> cbl<30> in1<13> in2<13> sl<61> vdd vss wl<13> / cell_PIM2
XI25192 vss vss in1<35> in2<35> vss vdd vss wl<35> / cell_PIM2
XI25191 vss vss in1<36> in2<36> vss vdd vss wl<36> / cell_PIM2
XI25190 vss vss in1<37> in2<37> vss vdd vss wl<37> / cell_PIM2
XI25189 vss vss in1<38> in2<38> vss vdd vss wl<38> / cell_PIM2
XI25193 vss vss in1<34> in2<34> vss vdd vss wl<34> / cell_PIM2
XI25188 vss vss in1<39> in2<39> vss vdd vss wl<39> / cell_PIM2
XI25187 vss vss in1<40> in2<40> vss vdd vss wl<40> / cell_PIM2
XI25186 vss vss in1<41> in2<41> vss vdd vss wl<41> / cell_PIM2
XI25185 vss vss in1<42> in2<42> vss vdd vss wl<42> / cell_PIM2
XI25184 vss vss in1<43> in2<43> vss vdd vss wl<43> / cell_PIM2
XI24533 bl<59> cbl<29> in1<14> in2<14> sl<59> vdd vss wl<14> / cell_PIM2
XI25182 vss vss in1<45> in2<45> vss vdd vss wl<45> / cell_PIM2
XI25181 vss vss in1<46> in2<46> vss vdd vss wl<46> / cell_PIM2
XI25180 vss vss in1<47> in2<47> vss vdd vss wl<47> / cell_PIM2
XI25179 vss vss in1<48> in2<48> vss vdd vss wl<48> / cell_PIM2
XI25183 vss vss in1<44> in2<44> vss vdd vss wl<44> / cell_PIM2
XI25177 vss vss in1<50> in2<50> vss vdd vss wl<50> / cell_PIM2
XI25176 vss vss in1<51> in2<51> vss vdd vss wl<51> / cell_PIM2
XI25175 vss vss in1<52> in2<52> vss vdd vss wl<52> / cell_PIM2
XI25174 vss vss in1<53> in2<53> vss vdd vss wl<53> / cell_PIM2
XI25178 vss vss in1<49> in2<49> vss vdd vss wl<49> / cell_PIM2
XI24523 bl<57> cbl<28> in1<14> in2<14> sl<57> vdd vss wl<14> / cell_PIM2
XI25172 vss vss in1<55> in2<55> vss vdd vss wl<55> / cell_PIM2
XI25171 vss vss in1<56> in2<56> vss vdd vss wl<56> / cell_PIM2
XI25170 vss vss in1<57> in2<57> vss vdd vss wl<57> / cell_PIM2
XI25169 vss vss in1<58> in2<58> vss vdd vss wl<58> / cell_PIM2
XI25173 vss vss in1<54> in2<54> vss vdd vss wl<54> / cell_PIM2
XI25168 vss vss in1<59> in2<59> vss vdd vss wl<59> / cell_PIM2
XI25167 vss vss in1<60> in2<60> vss vdd vss wl<60> / cell_PIM2
XI25166 vss vss in1<61> in2<61> vss vdd vss wl<61> / cell_PIM2
XI25165 vss vss in1<62> in2<62> vss vdd vss wl<62> / cell_PIM2
XI25164 vss vss in1<63> in2<63> vss vdd vss wl<63> / cell_PIM2
XI24513 bl<55> cbl<27> in1<14> in2<14> sl<55> vdd vss wl<14> / cell_PIM2
XI25162 vss vss in1<65> in2<65> vss vdd vss wl<65> / cell_PIM2
XI25161 vss vss in1<66> in2<66> vss vdd vss wl<66> / cell_PIM2
XI25160 vss vss in1<67> in2<67> vss vdd vss wl<67> / cell_PIM2
XI25159 vss vss in1<68> in2<68> vss vdd vss wl<68> / cell_PIM2
XI25163 vss vss in1<64> in2<64> vss vdd vss wl<64> / cell_PIM2
XI25157 vss vss in1<70> in2<70> vss vdd vss wl<70> / cell_PIM2
XI25156 vss vss in1<71> in2<71> vss vdd vss wl<71> / cell_PIM2
XI25155 vss vss in1<72> in2<72> vss vdd vss wl<72> / cell_PIM2
XI25154 vss vss in1<73> in2<73> vss vdd vss wl<73> / cell_PIM2
XI25158 vss vss in1<69> in2<69> vss vdd vss wl<69> / cell_PIM2
XI24503 bl<53> cbl<26> in1<13> in2<13> sl<53> vdd vss wl<13> / cell_PIM2
XI25152 vss vss in1<75> in2<75> vss vdd vss wl<75> / cell_PIM2
XI25151 vss vss in1<76> in2<76> vss vdd vss wl<76> / cell_PIM2
XI25150 vss vss in1<77> in2<77> vss vdd vss wl<77> / cell_PIM2
XI25149 vss vss in1<78> in2<78> vss vdd vss wl<78> / cell_PIM2
XI25153 vss vss in1<74> in2<74> vss vdd vss wl<74> / cell_PIM2
XI25148 vss vss in1<79> in2<79> vss vdd vss wl<79> / cell_PIM2
XI25147 vss vss in1<80> in2<80> vss vdd vss wl<80> / cell_PIM2
XI25146 vss vss in1<81> in2<81> vss vdd vss wl<81> / cell_PIM2
XI25145 vss vss in1<82> in2<82> vss vdd vss wl<82> / cell_PIM2
XI25144 vss vss in1<83> in2<83> vss vdd vss wl<83> / cell_PIM2
XI24493 bl<51> cbl<25> in1<14> in2<14> sl<51> vdd vss wl<14> / cell_PIM2
XI25142 vss vss in1<85> in2<85> vss vdd vss wl<85> / cell_PIM2
XI25141 vss vss in1<86> in2<86> vss vdd vss wl<86> / cell_PIM2
XI25140 vss vss in1<87> in2<87> vss vdd vss wl<87> / cell_PIM2
XI25139 vss vss in1<88> in2<88> vss vdd vss wl<88> / cell_PIM2
XI25143 vss vss in1<84> in2<84> vss vdd vss wl<84> / cell_PIM2
XI25137 vss vss in1<90> in2<90> vss vdd vss wl<90> / cell_PIM2
XI25136 vss vss in1<91> in2<91> vss vdd vss wl<91> / cell_PIM2
XI25135 vss vss in1<92> in2<92> vss vdd vss wl<92> / cell_PIM2
XI25134 vss vss in1<93> in2<93> vss vdd vss wl<93> / cell_PIM2
XI25138 vss vss in1<89> in2<89> vss vdd vss wl<89> / cell_PIM2
XI24483 bl<49> cbl<24> in1<13> in2<13> sl<49> vdd vss wl<13> / cell_PIM2
XI25132 vss vss in1<95> in2<95> vss vdd vss wl<95> / cell_PIM2
XI25131 vss vss in1<96> in2<96> vss vdd vss wl<96> / cell_PIM2
XI25130 vss vss in1<97> in2<97> vss vdd vss wl<97> / cell_PIM2
XI25129 vss vss in1<98> in2<98> vss vdd vss wl<98> / cell_PIM2
XI25133 vss vss in1<94> in2<94> vss vdd vss wl<94> / cell_PIM2
XI25128 vss vss in1<99> in2<99> vss vdd vss wl<99> / cell_PIM2
XI25127 vss vss in1<100> in2<100> vss vdd vss wl<100> / cell_PIM2
XI25126 vss vss in1<101> in2<101> vss vdd vss wl<101> / cell_PIM2
XI25125 vss vss in1<102> in2<102> vss vdd vss wl<102> / cell_PIM2
XI25124 vss vss in1<103> in2<103> vss vdd vss wl<103> / cell_PIM2
XI24473 bl<47> cbl<23> in1<14> in2<14> sl<47> vdd vss wl<14> / cell_PIM2
XI25122 vss vss in1<105> in2<105> vss vdd vss wl<105> / cell_PIM2
XI25121 vss vss in1<106> in2<106> vss vdd vss wl<106> / cell_PIM2
XI25120 vss vss in1<107> in2<107> vss vdd vss wl<107> / cell_PIM2
XI25119 vss vss in1<108> in2<108> vss vdd vss wl<108> / cell_PIM2
XI25123 vss vss in1<104> in2<104> vss vdd vss wl<104> / cell_PIM2
XI25117 vss vss in1<110> in2<110> vss vdd vss wl<110> / cell_PIM2
XI25116 vss vss in1<111> in2<111> vss vdd vss wl<111> / cell_PIM2
XI25115 vss vss in1<112> in2<112> vss vdd vss wl<112> / cell_PIM2
XI25114 vss vss in1<113> in2<113> vss vdd vss wl<113> / cell_PIM2
XI25118 vss vss in1<109> in2<109> vss vdd vss wl<109> / cell_PIM2
XI24463 bl<45> cbl<22> in1<13> in2<13> sl<45> vdd vss wl<13> / cell_PIM2
XI25112 vss vss in1<115> in2<115> vss vdd vss wl<115> / cell_PIM2
XI25111 vss vss in1<116> in2<116> vss vdd vss wl<116> / cell_PIM2
XI25110 vss vss in1<117> in2<117> vss vdd vss wl<117> / cell_PIM2
XI25109 vss vss in1<118> in2<118> vss vdd vss wl<118> / cell_PIM2
XI25113 vss vss in1<114> in2<114> vss vdd vss wl<114> / cell_PIM2
XI25108 vss vss in1<119> in2<119> vss vdd vss wl<119> / cell_PIM2
XI25107 vss vss in1<120> in2<120> vss vdd vss wl<120> / cell_PIM2
XI25106 vss vss in1<121> in2<121> vss vdd vss wl<121> / cell_PIM2
XI25105 vss vss in1<122> in2<122> vss vdd vss wl<122> / cell_PIM2
XI25104 vss vss in1<123> in2<123> vss vdd vss wl<123> / cell_PIM2
XI24453 bl<43> cbl<21> in1<14> in2<14> sl<43> vdd vss wl<14> / cell_PIM2
XI25102 vss vss in1<127> in2<127> vss vdd vss wl<127> / cell_PIM2
XI25101 vss vss in1<126> in2<126> vss vdd vss wl<126> / cell_PIM2
XI25100 vss vss in1<125> in2<125> vss vdd vss wl<125> / cell_PIM2
XI25099 vss vss in1<124> in2<124> vss vdd vss wl<124> / cell_PIM2
XI25103 vss vss vdd vdd vss vdd vss vss / cell_PIM2
XI25096 bl<61> cbl<30> vdd vdd sl<61> vdd vss vss / cell_PIM2
XI25094 bl<59> cbl<29> vdd vdd sl<59> vdd vss vss / cell_PIM2
XI25098 bl<63> cbl<31> vdd vdd sl<63> vdd vss vss / cell_PIM2
XI24443 bl<41> cbl<20> in1<14> in2<14> sl<41> vdd vss wl<14> / cell_PIM2
XI25092 bl<57> cbl<28> vdd vdd sl<57> vdd vss vss / cell_PIM2
XI25090 bl<55> cbl<27> vdd vdd sl<55> vdd vss vss / cell_PIM2
XI25088 bl<53> cbl<26> vdd vdd sl<53> vdd vss vss / cell_PIM2
XI25086 bl<51> cbl<25> vdd vdd sl<51> vdd vss vss / cell_PIM2
XI25084 bl<49> cbl<24> vdd vdd sl<49> vdd vss vss / cell_PIM2
XI24433 bl<39> cbl<19> in1<14> in2<14> sl<39> vdd vss wl<14> / cell_PIM2
XI25082 bl<47> cbl<23> vdd vdd sl<47> vdd vss vss / cell_PIM2
XI25080 bl<45> cbl<22> vdd vdd sl<45> vdd vss vss / cell_PIM2
XI25076 bl<41> cbl<20> vdd vdd sl<41> vdd vss vss / cell_PIM2
XI25074 bl<39> cbl<19> vdd vdd sl<39> vdd vss vss / cell_PIM2
XI25078 bl<43> cbl<21> vdd vdd sl<43> vdd vss vss / cell_PIM2
XI24423 bl<37> cbl<18> in1<13> in2<13> sl<37> vdd vss wl<13> / cell_PIM2
XI25072 bl<37> cbl<18> vdd vdd sl<37> vdd vss vss / cell_PIM2
XI25070 bl<35> cbl<17> vdd vdd sl<35> vdd vss vss / cell_PIM2
XI25068 bl<33> cbl<16> vdd vdd sl<33> vdd vss vss / cell_PIM2
XI25066 bl<31> cbl<15> vdd vdd sl<31> vdd vss vss / cell_PIM2
XI25064 bl<29> cbl<14> vdd vdd sl<29> vdd vss vss / cell_PIM2
XI24413 bl<35> cbl<17> in1<14> in2<14> sl<35> vdd vss wl<14> / cell_PIM2
XI25062 bl<27> cbl<13> vdd vdd sl<27> vdd vss vss / cell_PIM2
XI25060 bl<25> cbl<12> vdd vdd sl<25> vdd vss vss / cell_PIM2
XI25056 bl<21> cbl<10> vdd vdd sl<21> vdd vss vss / cell_PIM2
XI25054 bl<19> cbl<9> vdd vdd sl<19> vdd vss vss / cell_PIM2
XI25058 bl<23> cbl<11> vdd vdd sl<23> vdd vss vss / cell_PIM2
XI24403 bl<33> cbl<16> in1<13> in2<13> sl<33> vdd vss wl<13> / cell_PIM2
XI25052 bl<17> cbl<8> vdd vdd sl<17> vdd vss vss / cell_PIM2
XI25050 bl<15> cbl<7> vdd vdd sl<15> vdd vss vss / cell_PIM2
XI25048 bl<13> cbl<6> vdd vdd sl<13> vdd vss vss / cell_PIM2
XI25046 bl<11> cbl<5> vdd vdd sl<11> vdd vss vss / cell_PIM2
XI25044 bl<9> cbl<4> vdd vdd sl<9> vdd vss vss / cell_PIM2
XI24393 bl<63> cbl<31> in1<19> in2<19> sl<63> vdd vss wl<19> / cell_PIM2
XI25042 bl<7> cbl<3> vdd vdd sl<7> vdd vss vss / cell_PIM2
XI25040 bl<5> cbl<2> vdd vdd sl<5> vdd vss vss / cell_PIM2
XI25036 bl<1> cbl<0> vdd vdd sl<1> vdd vss vss / cell_PIM2
XI25034 bl<63> cbl<31> vdd vdd sl<63> vdd vss vss / cell_PIM2
XI25038 bl<3> cbl<1> vdd vdd sl<3> vdd vss vss / cell_PIM2
XI23404 bl<45> cbl<22> in1<48> in2<48> sl<45> vdd vss wl<48> / cell_PIM2
XI24053 bl<53> cbl<26> in1<30> in2<30> sl<53> vdd vss wl<30> / cell_PIM2
XI24052 bl<53> cbl<26> in1<29> in2<29> sl<53> vdd vss wl<29> / cell_PIM2
XI24702 bl<61> cbl<30> in1<12> in2<12> sl<61> vdd vss wl<12> / cell_PIM2
XI24701 bl<61> cbl<30> in1<11> in2<11> sl<61> vdd vss wl<11> / cell_PIM2
XI24700 bl<61> cbl<30> in1<10> in2<10> sl<61> vdd vss wl<10> / cell_PIM2
XI24694 bl<59> cbl<29> in1<8> in2<8> sl<59> vdd vss wl<8> / cell_PIM2
XI24046 bl<51> cbl<25> in1<27> in2<27> sl<51> vdd vss wl<27> / cell_PIM2
XI24045 bl<51> cbl<25> in1<28> in2<28> sl<51> vdd vss wl<28> / cell_PIM2
XI24044 bl<51> cbl<25> in1<29> in2<29> sl<51> vdd vss wl<29> / cell_PIM2
XI23398 bl<43> cbl<21> in1<46> in2<46> sl<43> vdd vss wl<46> / cell_PIM2
XI23397 bl<43> cbl<21> in1<47> in2<47> sl<43> vdd vss wl<47> / cell_PIM2
XI22878 bl<61> cbl<30> in1<65> in2<65> sl<61> vdd vss wl<65> / cell_PIM2
XI23396 bl<43> cbl<21> in1<48> in2<48> sl<43> vdd vss wl<48> / cell_PIM2
XI23395 bl<43> cbl<21> in1<49> in2<49> sl<43> vdd vss wl<49> / cell_PIM2
XI23394 bl<43> cbl<21> in1<50> in2<50> sl<43> vdd vss wl<50> / cell_PIM2
XI24043 bl<51> cbl<25> in1<30> in2<30> sl<51> vdd vss wl<30> / cell_PIM2
XI24042 bl<51> cbl<25> in1<31> in2<31> sl<51> vdd vss wl<31> / cell_PIM2
XI24692 bl<59> cbl<29> in1<10> in2<10> sl<59> vdd vss wl<10> / cell_PIM2
XI24691 bl<59> cbl<29> in1<11> in2<11> sl<59> vdd vss wl<11> / cell_PIM2
XI24690 bl<59> cbl<29> in1<12> in2<12> sl<59> vdd vss wl<12> / cell_PIM2
XI22868 bl<59> cbl<29> in1<67> in2<67> sl<59> vdd vss wl<67> / cell_PIM2
XI24036 bl<49> cbl<24> in1<28> in2<28> sl<49> vdd vss wl<28> / cell_PIM2
XI24035 bl<49> cbl<24> in1<27> in2<27> sl<49> vdd vss wl<27> / cell_PIM2
XI24034 bl<49> cbl<24> in1<31> in2<31> sl<49> vdd vss wl<31> / cell_PIM2
XI24684 bl<57> cbl<28> in1<8> in2<8> sl<57> vdd vss wl<8> / cell_PIM2
XI23388 bl<41> cbl<20> in1<46> in2<46> sl<41> vdd vss wl<46> / cell_PIM2
XI23387 bl<41> cbl<20> in1<47> in2<47> sl<41> vdd vss wl<47> / cell_PIM2
XI23386 bl<41> cbl<20> in1<48> in2<48> sl<41> vdd vss wl<48> / cell_PIM2
XI23385 bl<41> cbl<20> in1<49> in2<49> sl<41> vdd vss wl<49> / cell_PIM2
XI24033 bl<49> cbl<24> in1<30> in2<30> sl<49> vdd vss wl<30> / cell_PIM2
XI24032 bl<49> cbl<24> in1<29> in2<29> sl<49> vdd vss wl<29> / cell_PIM2
XI24682 bl<57> cbl<28> in1<10> in2<10> sl<57> vdd vss wl<10> / cell_PIM2
XI24681 bl<57> cbl<28> in1<11> in2<11> sl<57> vdd vss wl<11> / cell_PIM2
XI24680 bl<57> cbl<28> in1<12> in2<12> sl<57> vdd vss wl<12> / cell_PIM2
XI24674 bl<55> cbl<27> in1<8> in2<8> sl<55> vdd vss wl<8> / cell_PIM2
XI24026 bl<47> cbl<23> in1<27> in2<27> sl<47> vdd vss wl<27> / cell_PIM2
XI24025 bl<47> cbl<23> in1<28> in2<28> sl<47> vdd vss wl<28> / cell_PIM2
XI24024 bl<47> cbl<23> in1<29> in2<29> sl<47> vdd vss wl<29> / cell_PIM2
XI23384 bl<41> cbl<20> in1<50> in2<50> sl<41> vdd vss wl<50> / cell_PIM2
XI22858 bl<57> cbl<28> in1<67> in2<67> sl<57> vdd vss wl<67> / cell_PIM2
XI23378 bl<39> cbl<19> in1<46> in2<46> sl<39> vdd vss wl<46> / cell_PIM2
XI23377 bl<39> cbl<19> in1<47> in2<47> sl<39> vdd vss wl<47> / cell_PIM2
XI24023 bl<47> cbl<23> in1<30> in2<30> sl<47> vdd vss wl<30> / cell_PIM2
XI24022 bl<47> cbl<23> in1<31> in2<31> sl<47> vdd vss wl<31> / cell_PIM2
XI24672 bl<55> cbl<27> in1<10> in2<10> sl<55> vdd vss wl<10> / cell_PIM2
XI24671 bl<55> cbl<27> in1<11> in2<11> sl<55> vdd vss wl<11> / cell_PIM2
XI24670 bl<55> cbl<27> in1<12> in2<12> sl<55> vdd vss wl<12> / cell_PIM2
XI22848 bl<55> cbl<27> in1<67> in2<67> sl<55> vdd vss wl<67> / cell_PIM2
XI23376 bl<39> cbl<19> in1<48> in2<48> sl<39> vdd vss wl<48> / cell_PIM2
XI23375 bl<39> cbl<19> in1<49> in2<49> sl<39> vdd vss wl<49> / cell_PIM2
XI23374 bl<39> cbl<19> in1<50> in2<50> sl<39> vdd vss wl<50> / cell_PIM2
XI24016 bl<45> cbl<22> in1<28> in2<28> sl<45> vdd vss wl<28> / cell_PIM2
XI24015 bl<45> cbl<22> in1<27> in2<27> sl<45> vdd vss wl<27> / cell_PIM2
XI24014 bl<45> cbl<22> in1<31> in2<31> sl<45> vdd vss wl<31> / cell_PIM2
XI24664 bl<53> cbl<26> in1<9> in2<9> sl<53> vdd vss wl<9> / cell_PIM2
XI24013 bl<45> cbl<22> in1<30> in2<30> sl<45> vdd vss wl<30> / cell_PIM2
XI24012 bl<45> cbl<22> in1<29> in2<29> sl<45> vdd vss wl<29> / cell_PIM2
XI24662 bl<53> cbl<26> in1<12> in2<12> sl<53> vdd vss wl<12> / cell_PIM2
XI24661 bl<53> cbl<26> in1<11> in2<11> sl<53> vdd vss wl<11> / cell_PIM2
XI24660 bl<53> cbl<26> in1<10> in2<10> sl<53> vdd vss wl<10> / cell_PIM2
XI24654 bl<51> cbl<25> in1<8> in2<8> sl<51> vdd vss wl<8> / cell_PIM2
XI24006 bl<43> cbl<21> in1<27> in2<27> sl<43> vdd vss wl<27> / cell_PIM2
XI24005 bl<43> cbl<21> in1<28> in2<28> sl<43> vdd vss wl<28> / cell_PIM2
XI24004 bl<43> cbl<21> in1<29> in2<29> sl<43> vdd vss wl<29> / cell_PIM2
XI23368 bl<37> cbl<18> in1<47> in2<47> sl<37> vdd vss wl<47> / cell_PIM2
XI23367 bl<37> cbl<18> in1<46> in2<46> sl<37> vdd vss wl<46> / cell_PIM2
XI23366 bl<37> cbl<18> in1<50> in2<50> sl<37> vdd vss wl<50> / cell_PIM2
XI23365 bl<37> cbl<18> in1<49> in2<49> sl<37> vdd vss wl<49> / cell_PIM2
XI22838 bl<53> cbl<26> in1<65> in2<65> sl<53> vdd vss wl<65> / cell_PIM2
XI23364 bl<37> cbl<18> in1<48> in2<48> sl<37> vdd vss wl<48> / cell_PIM2
XI24003 bl<43> cbl<21> in1<30> in2<30> sl<43> vdd vss wl<30> / cell_PIM2
XI24002 bl<43> cbl<21> in1<31> in2<31> sl<43> vdd vss wl<31> / cell_PIM2
XI24652 bl<51> cbl<25> in1<10> in2<10> sl<51> vdd vss wl<10> / cell_PIM2
XI24651 bl<51> cbl<25> in1<11> in2<11> sl<51> vdd vss wl<11> / cell_PIM2
XI24650 bl<51> cbl<25> in1<12> in2<12> sl<51> vdd vss wl<12> / cell_PIM2
XI22828 bl<51> cbl<25> in1<67> in2<67> sl<51> vdd vss wl<67> / cell_PIM2
XI23358 bl<35> cbl<17> in1<46> in2<46> sl<35> vdd vss wl<46> / cell_PIM2
XI23357 bl<35> cbl<17> in1<47> in2<47> sl<35> vdd vss wl<47> / cell_PIM2
XI23996 bl<41> cbl<20> in1<27> in2<27> sl<41> vdd vss wl<27> / cell_PIM2
XI23995 bl<41> cbl<20> in1<28> in2<28> sl<41> vdd vss wl<28> / cell_PIM2
XI23994 bl<41> cbl<20> in1<29> in2<29> sl<41> vdd vss wl<29> / cell_PIM2
XI24644 bl<49> cbl<24> in1<9> in2<9> sl<49> vdd vss wl<9> / cell_PIM2
XI23356 bl<35> cbl<17> in1<48> in2<48> sl<35> vdd vss wl<48> / cell_PIM2
XI23355 bl<35> cbl<17> in1<49> in2<49> sl<35> vdd vss wl<49> / cell_PIM2
XI23354 bl<35> cbl<17> in1<50> in2<50> sl<35> vdd vss wl<50> / cell_PIM2
XI23993 bl<41> cbl<20> in1<30> in2<30> sl<41> vdd vss wl<30> / cell_PIM2
XI23992 bl<41> cbl<20> in1<31> in2<31> sl<41> vdd vss wl<31> / cell_PIM2
XI24642 bl<49> cbl<24> in1<12> in2<12> sl<49> vdd vss wl<12> / cell_PIM2
XI24641 bl<49> cbl<24> in1<11> in2<11> sl<49> vdd vss wl<11> / cell_PIM2
XI24640 bl<49> cbl<24> in1<10> in2<10> sl<49> vdd vss wl<10> / cell_PIM2
XI24634 bl<47> cbl<23> in1<8> in2<8> sl<47> vdd vss wl<8> / cell_PIM2
XI23986 bl<39> cbl<19> in1<27> in2<27> sl<39> vdd vss wl<27> / cell_PIM2
XI23985 bl<39> cbl<19> in1<28> in2<28> sl<39> vdd vss wl<28> / cell_PIM2
XI23984 bl<39> cbl<19> in1<29> in2<29> sl<39> vdd vss wl<29> / cell_PIM2
XI22818 bl<49> cbl<24> in1<65> in2<65> sl<49> vdd vss wl<65> / cell_PIM2
XI23348 bl<33> cbl<16> in1<47> in2<47> sl<33> vdd vss wl<47> / cell_PIM2
XI23347 bl<33> cbl<16> in1<46> in2<46> sl<33> vdd vss wl<46> / cell_PIM2
XI23346 bl<33> cbl<16> in1<50> in2<50> sl<33> vdd vss wl<50> / cell_PIM2
XI23345 bl<33> cbl<16> in1<49> in2<49> sl<33> vdd vss wl<49> / cell_PIM2
XI23983 bl<39> cbl<19> in1<30> in2<30> sl<39> vdd vss wl<30> / cell_PIM2
XI23982 bl<39> cbl<19> in1<31> in2<31> sl<39> vdd vss wl<31> / cell_PIM2
XI24632 bl<47> cbl<23> in1<10> in2<10> sl<47> vdd vss wl<10> / cell_PIM2
XI24631 bl<47> cbl<23> in1<11> in2<11> sl<47> vdd vss wl<11> / cell_PIM2
XI24630 bl<47> cbl<23> in1<12> in2<12> sl<47> vdd vss wl<12> / cell_PIM2
XI22808 bl<47> cbl<23> in1<67> in2<67> sl<47> vdd vss wl<67> / cell_PIM2
XI23344 bl<33> cbl<16> in1<48> in2<48> sl<33> vdd vss wl<48> / cell_PIM2
XI23976 bl<37> cbl<18> in1<28> in2<28> sl<37> vdd vss wl<28> / cell_PIM2
XI23975 bl<37> cbl<18> in1<27> in2<27> sl<37> vdd vss wl<27> / cell_PIM2
XI23974 bl<37> cbl<18> in1<31> in2<31> sl<37> vdd vss wl<31> / cell_PIM2
XI24624 bl<45> cbl<22> in1<9> in2<9> sl<45> vdd vss wl<9> / cell_PIM2
XI23338 bl<63> cbl<31> in1<51> in2<51> sl<63> vdd vss wl<51> / cell_PIM2
XI23337 bl<63> cbl<31> in1<52> in2<52> sl<63> vdd vss wl<52> / cell_PIM2
XI23973 bl<37> cbl<18> in1<30> in2<30> sl<37> vdd vss wl<30> / cell_PIM2
XI23972 bl<37> cbl<18> in1<29> in2<29> sl<37> vdd vss wl<29> / cell_PIM2
XI24622 bl<45> cbl<22> in1<12> in2<12> sl<45> vdd vss wl<12> / cell_PIM2
XI24621 bl<45> cbl<22> in1<11> in2<11> sl<45> vdd vss wl<11> / cell_PIM2
XI24620 bl<45> cbl<22> in1<10> in2<10> sl<45> vdd vss wl<10> / cell_PIM2
XI24614 bl<43> cbl<21> in1<8> in2<8> sl<43> vdd vss wl<8> / cell_PIM2
XI23966 bl<35> cbl<17> in1<27> in2<27> sl<35> vdd vss wl<27> / cell_PIM2
XI23965 bl<35> cbl<17> in1<28> in2<28> sl<35> vdd vss wl<28> / cell_PIM2
XI23964 bl<35> cbl<17> in1<29> in2<29> sl<35> vdd vss wl<29> / cell_PIM2
XI23336 bl<63> cbl<31> in1<53> in2<53> sl<63> vdd vss wl<53> / cell_PIM2
XI23335 bl<63> cbl<31> in1<54> in2<54> sl<63> vdd vss wl<54> / cell_PIM2
XI23334 bl<63> cbl<31> in1<55> in2<55> sl<63> vdd vss wl<55> / cell_PIM2
XI22798 bl<45> cbl<22> in1<65> in2<65> sl<45> vdd vss wl<65> / cell_PIM2
XI23963 bl<35> cbl<17> in1<30> in2<30> sl<35> vdd vss wl<30> / cell_PIM2
XI23962 bl<35> cbl<17> in1<31> in2<31> sl<35> vdd vss wl<31> / cell_PIM2
XI24612 bl<43> cbl<21> in1<10> in2<10> sl<43> vdd vss wl<10> / cell_PIM2
XI24611 bl<43> cbl<21> in1<11> in2<11> sl<43> vdd vss wl<11> / cell_PIM2
XI24610 bl<43> cbl<21> in1<12> in2<12> sl<43> vdd vss wl<12> / cell_PIM2
XI22788 bl<43> cbl<21> in1<67> in2<67> sl<43> vdd vss wl<67> / cell_PIM2
XI23328 bl<61> cbl<30> in1<52> in2<52> sl<61> vdd vss wl<52> / cell_PIM2
XI23327 bl<61> cbl<30> in1<51> in2<51> sl<61> vdd vss wl<51> / cell_PIM2
XI23326 bl<61> cbl<30> in1<55> in2<55> sl<61> vdd vss wl<55> / cell_PIM2
XI23325 bl<61> cbl<30> in1<54> in2<54> sl<61> vdd vss wl<54> / cell_PIM2
XI23956 bl<33> cbl<16> in1<28> in2<28> sl<33> vdd vss wl<28> / cell_PIM2
XI23955 bl<33> cbl<16> in1<27> in2<27> sl<33> vdd vss wl<27> / cell_PIM2
XI23954 bl<33> cbl<16> in1<31> in2<31> sl<33> vdd vss wl<31> / cell_PIM2
XI24604 bl<41> cbl<20> in1<8> in2<8> sl<41> vdd vss wl<8> / cell_PIM2
XI23324 bl<61> cbl<30> in1<53> in2<53> sl<61> vdd vss wl<53> / cell_PIM2
XI23953 bl<33> cbl<16> in1<30> in2<30> sl<33> vdd vss wl<30> / cell_PIM2
XI23952 bl<33> cbl<16> in1<29> in2<29> sl<33> vdd vss wl<29> / cell_PIM2
XI24602 bl<41> cbl<20> in1<10> in2<10> sl<41> vdd vss wl<10> / cell_PIM2
XI24601 bl<41> cbl<20> in1<11> in2<11> sl<41> vdd vss wl<11> / cell_PIM2
XI24600 bl<41> cbl<20> in1<12> in2<12> sl<41> vdd vss wl<12> / cell_PIM2
XI24594 bl<39> cbl<19> in1<8> in2<8> sl<39> vdd vss wl<8> / cell_PIM2
XI23946 bl<63> cbl<31> in1<32> in2<32> sl<63> vdd vss wl<32> / cell_PIM2
XI23945 bl<63> cbl<31> in1<33> in2<33> sl<63> vdd vss wl<33> / cell_PIM2
XI23944 bl<63> cbl<31> in1<34> in2<34> sl<63> vdd vss wl<34> / cell_PIM2
XI23318 bl<59> cbl<29> in1<51> in2<51> sl<59> vdd vss wl<51> / cell_PIM2
XI23317 bl<59> cbl<29> in1<52> in2<52> sl<59> vdd vss wl<52> / cell_PIM2
XI22778 bl<41> cbl<20> in1<67> in2<67> sl<41> vdd vss wl<67> / cell_PIM2
XI23316 bl<59> cbl<29> in1<53> in2<53> sl<59> vdd vss wl<53> / cell_PIM2
XI23315 bl<59> cbl<29> in1<54> in2<54> sl<59> vdd vss wl<54> / cell_PIM2
XI23314 bl<59> cbl<29> in1<55> in2<55> sl<59> vdd vss wl<55> / cell_PIM2
XI23943 bl<63> cbl<31> in1<35> in2<35> sl<63> vdd vss wl<35> / cell_PIM2
XI23942 bl<63> cbl<31> in1<36> in2<36> sl<63> vdd vss wl<36> / cell_PIM2
XI24592 bl<39> cbl<19> in1<10> in2<10> sl<39> vdd vss wl<10> / cell_PIM2
XI24591 bl<39> cbl<19> in1<11> in2<11> sl<39> vdd vss wl<11> / cell_PIM2
XI24590 bl<39> cbl<19> in1<12> in2<12> sl<39> vdd vss wl<12> / cell_PIM2
XI22768 bl<39> cbl<19> in1<67> in2<67> sl<39> vdd vss wl<67> / cell_PIM2
XI23936 bl<61> cbl<30> in1<33> in2<33> sl<61> vdd vss wl<33> / cell_PIM2
XI23935 bl<61> cbl<30> in1<32> in2<32> sl<61> vdd vss wl<32> / cell_PIM2
XI23934 bl<61> cbl<30> in1<36> in2<36> sl<61> vdd vss wl<36> / cell_PIM2
XI24584 bl<37> cbl<18> in1<9> in2<9> sl<37> vdd vss wl<9> / cell_PIM2
XI23308 bl<57> cbl<28> in1<51> in2<51> sl<57> vdd vss wl<51> / cell_PIM2
XI23307 bl<57> cbl<28> in1<52> in2<52> sl<57> vdd vss wl<52> / cell_PIM2
XI23306 bl<57> cbl<28> in1<53> in2<53> sl<57> vdd vss wl<53> / cell_PIM2
XI23305 bl<57> cbl<28> in1<54> in2<54> sl<57> vdd vss wl<54> / cell_PIM2
XI23933 bl<61> cbl<30> in1<35> in2<35> sl<61> vdd vss wl<35> / cell_PIM2
XI23932 bl<61> cbl<30> in1<34> in2<34> sl<61> vdd vss wl<34> / cell_PIM2
XI24582 bl<37> cbl<18> in1<12> in2<12> sl<37> vdd vss wl<12> / cell_PIM2
XI24581 bl<37> cbl<18> in1<11> in2<11> sl<37> vdd vss wl<11> / cell_PIM2
XI24580 bl<37> cbl<18> in1<10> in2<10> sl<37> vdd vss wl<10> / cell_PIM2
XI24574 bl<35> cbl<17> in1<8> in2<8> sl<35> vdd vss wl<8> / cell_PIM2
XI23926 bl<59> cbl<29> in1<32> in2<32> sl<59> vdd vss wl<32> / cell_PIM2
XI23925 bl<59> cbl<29> in1<33> in2<33> sl<59> vdd vss wl<33> / cell_PIM2
XI23924 bl<59> cbl<29> in1<34> in2<34> sl<59> vdd vss wl<34> / cell_PIM2
XI23304 bl<57> cbl<28> in1<55> in2<55> sl<57> vdd vss wl<55> / cell_PIM2
XI22758 bl<37> cbl<18> in1<65> in2<65> sl<37> vdd vss wl<65> / cell_PIM2
XI23298 bl<55> cbl<27> in1<51> in2<51> sl<55> vdd vss wl<51> / cell_PIM2
XI23297 bl<55> cbl<27> in1<52> in2<52> sl<55> vdd vss wl<52> / cell_PIM2
XI23923 bl<59> cbl<29> in1<35> in2<35> sl<59> vdd vss wl<35> / cell_PIM2
XI23922 bl<59> cbl<29> in1<36> in2<36> sl<59> vdd vss wl<36> / cell_PIM2
XI24572 bl<35> cbl<17> in1<10> in2<10> sl<35> vdd vss wl<10> / cell_PIM2
XI24571 bl<35> cbl<17> in1<11> in2<11> sl<35> vdd vss wl<11> / cell_PIM2
XI24570 bl<35> cbl<17> in1<12> in2<12> sl<35> vdd vss wl<12> / cell_PIM2
XI22748 bl<35> cbl<17> in1<67> in2<67> sl<35> vdd vss wl<67> / cell_PIM2
XI23296 bl<55> cbl<27> in1<53> in2<53> sl<55> vdd vss wl<53> / cell_PIM2
XI23295 bl<55> cbl<27> in1<54> in2<54> sl<55> vdd vss wl<54> / cell_PIM2
XI23294 bl<55> cbl<27> in1<55> in2<55> sl<55> vdd vss wl<55> / cell_PIM2
XI23916 bl<57> cbl<28> in1<32> in2<32> sl<57> vdd vss wl<32> / cell_PIM2
XI23915 bl<57> cbl<28> in1<33> in2<33> sl<57> vdd vss wl<33> / cell_PIM2
XI23914 bl<57> cbl<28> in1<34> in2<34> sl<57> vdd vss wl<34> / cell_PIM2
XI24564 bl<33> cbl<16> in1<9> in2<9> sl<33> vdd vss wl<9> / cell_PIM2
XI23913 bl<57> cbl<28> in1<35> in2<35> sl<57> vdd vss wl<35> / cell_PIM2
XI23912 bl<57> cbl<28> in1<36> in2<36> sl<57> vdd vss wl<36> / cell_PIM2
XI24562 bl<33> cbl<16> in1<12> in2<12> sl<33> vdd vss wl<12> / cell_PIM2
XI24561 bl<33> cbl<16> in1<11> in2<11> sl<33> vdd vss wl<11> / cell_PIM2
XI24560 bl<33> cbl<16> in1<10> in2<10> sl<33> vdd vss wl<10> / cell_PIM2
XI24554 bl<63> cbl<31> in1<13> in2<13> sl<63> vdd vss wl<13> / cell_PIM2
XI23906 bl<55> cbl<27> in1<32> in2<32> sl<55> vdd vss wl<32> / cell_PIM2
XI23905 bl<55> cbl<27> in1<33> in2<33> sl<55> vdd vss wl<33> / cell_PIM2
XI23904 bl<55> cbl<27> in1<34> in2<34> sl<55> vdd vss wl<34> / cell_PIM2
XI23288 bl<53> cbl<26> in1<52> in2<52> sl<53> vdd vss wl<52> / cell_PIM2
XI23287 bl<53> cbl<26> in1<51> in2<51> sl<53> vdd vss wl<51> / cell_PIM2
XI23286 bl<53> cbl<26> in1<55> in2<55> sl<53> vdd vss wl<55> / cell_PIM2
XI23285 bl<53> cbl<26> in1<54> in2<54> sl<53> vdd vss wl<54> / cell_PIM2
XI22738 bl<33> cbl<16> in1<65> in2<65> sl<33> vdd vss wl<65> / cell_PIM2
XI23284 bl<53> cbl<26> in1<53> in2<53> sl<53> vdd vss wl<53> / cell_PIM2
XI23903 bl<55> cbl<27> in1<35> in2<35> sl<55> vdd vss wl<35> / cell_PIM2
XI23902 bl<55> cbl<27> in1<36> in2<36> sl<55> vdd vss wl<36> / cell_PIM2
XI24552 bl<63> cbl<31> in1<15> in2<15> sl<63> vdd vss wl<15> / cell_PIM2
XI24551 bl<63> cbl<31> in1<16> in2<16> sl<63> vdd vss wl<16> / cell_PIM2
XI24550 bl<63> cbl<31> in1<17> in2<17> sl<63> vdd vss wl<17> / cell_PIM2
XI22728 bl<63> cbl<31> in1<72> in2<72> sl<63> vdd vss wl<72> / cell_PIM2
XI23278 bl<51> cbl<25> in1<51> in2<51> sl<51> vdd vss wl<51> / cell_PIM2
XI23277 bl<51> cbl<25> in1<52> in2<52> sl<51> vdd vss wl<52> / cell_PIM2
XI23896 bl<53> cbl<26> in1<33> in2<33> sl<53> vdd vss wl<33> / cell_PIM2
XI23895 bl<53> cbl<26> in1<32> in2<32> sl<53> vdd vss wl<32> / cell_PIM2
XI23894 bl<53> cbl<26> in1<36> in2<36> sl<53> vdd vss wl<36> / cell_PIM2
XI24544 bl<61> cbl<30> in1<14> in2<14> sl<61> vdd vss wl<14> / cell_PIM2
XI23276 bl<51> cbl<25> in1<53> in2<53> sl<51> vdd vss wl<53> / cell_PIM2
XI23275 bl<51> cbl<25> in1<54> in2<54> sl<51> vdd vss wl<54> / cell_PIM2
XI23274 bl<51> cbl<25> in1<55> in2<55> sl<51> vdd vss wl<55> / cell_PIM2
XI23893 bl<53> cbl<26> in1<35> in2<35> sl<53> vdd vss wl<35> / cell_PIM2
XI23892 bl<53> cbl<26> in1<34> in2<34> sl<53> vdd vss wl<34> / cell_PIM2
XI24542 bl<61> cbl<30> in1<17> in2<17> sl<61> vdd vss wl<17> / cell_PIM2
XI24541 bl<61> cbl<30> in1<16> in2<16> sl<61> vdd vss wl<16> / cell_PIM2
XI24540 bl<61> cbl<30> in1<15> in2<15> sl<61> vdd vss wl<15> / cell_PIM2
XI24534 bl<59> cbl<29> in1<13> in2<13> sl<59> vdd vss wl<13> / cell_PIM2
XI23886 bl<51> cbl<25> in1<32> in2<32> sl<51> vdd vss wl<32> / cell_PIM2
XI23885 bl<51> cbl<25> in1<33> in2<33> sl<51> vdd vss wl<33> / cell_PIM2
XI23884 bl<51> cbl<25> in1<34> in2<34> sl<51> vdd vss wl<34> / cell_PIM2
XI22718 bl<61> cbl<30> in1<74> in2<74> sl<61> vdd vss wl<74> / cell_PIM2
XI23268 bl<49> cbl<24> in1<52> in2<52> sl<49> vdd vss wl<52> / cell_PIM2
XI23267 bl<49> cbl<24> in1<51> in2<51> sl<49> vdd vss wl<51> / cell_PIM2
XI23266 bl<49> cbl<24> in1<55> in2<55> sl<49> vdd vss wl<55> / cell_PIM2
XI23265 bl<49> cbl<24> in1<54> in2<54> sl<49> vdd vss wl<54> / cell_PIM2
XI23883 bl<51> cbl<25> in1<35> in2<35> sl<51> vdd vss wl<35> / cell_PIM2
XI23882 bl<51> cbl<25> in1<36> in2<36> sl<51> vdd vss wl<36> / cell_PIM2
XI24532 bl<59> cbl<29> in1<15> in2<15> sl<59> vdd vss wl<15> / cell_PIM2
XI24531 bl<59> cbl<29> in1<16> in2<16> sl<59> vdd vss wl<16> / cell_PIM2
XI24530 bl<59> cbl<29> in1<17> in2<17> sl<59> vdd vss wl<17> / cell_PIM2
XI22708 bl<59> cbl<29> in1<72> in2<72> sl<59> vdd vss wl<72> / cell_PIM2
XI23264 bl<49> cbl<24> in1<53> in2<53> sl<49> vdd vss wl<53> / cell_PIM2
XI23876 bl<49> cbl<24> in1<33> in2<33> sl<49> vdd vss wl<33> / cell_PIM2
XI23875 bl<49> cbl<24> in1<32> in2<32> sl<49> vdd vss wl<32> / cell_PIM2
XI23874 bl<49> cbl<24> in1<36> in2<36> sl<49> vdd vss wl<36> / cell_PIM2
XI24524 bl<57> cbl<28> in1<13> in2<13> sl<57> vdd vss wl<13> / cell_PIM2
XI23258 bl<47> cbl<23> in1<51> in2<51> sl<47> vdd vss wl<51> / cell_PIM2
XI23257 bl<47> cbl<23> in1<52> in2<52> sl<47> vdd vss wl<52> / cell_PIM2
XI23873 bl<49> cbl<24> in1<35> in2<35> sl<49> vdd vss wl<35> / cell_PIM2
XI23872 bl<49> cbl<24> in1<34> in2<34> sl<49> vdd vss wl<34> / cell_PIM2
XI24522 bl<57> cbl<28> in1<15> in2<15> sl<57> vdd vss wl<15> / cell_PIM2
XI24521 bl<57> cbl<28> in1<16> in2<16> sl<57> vdd vss wl<16> / cell_PIM2
XI24520 bl<57> cbl<28> in1<17> in2<17> sl<57> vdd vss wl<17> / cell_PIM2
XI24514 bl<55> cbl<27> in1<13> in2<13> sl<55> vdd vss wl<13> / cell_PIM2
XI23866 bl<47> cbl<23> in1<32> in2<32> sl<47> vdd vss wl<32> / cell_PIM2
XI23865 bl<47> cbl<23> in1<33> in2<33> sl<47> vdd vss wl<33> / cell_PIM2
XI23864 bl<47> cbl<23> in1<34> in2<34> sl<47> vdd vss wl<34> / cell_PIM2
XI23256 bl<47> cbl<23> in1<53> in2<53> sl<47> vdd vss wl<53> / cell_PIM2
XI23255 bl<47> cbl<23> in1<54> in2<54> sl<47> vdd vss wl<54> / cell_PIM2
XI23254 bl<47> cbl<23> in1<55> in2<55> sl<47> vdd vss wl<55> / cell_PIM2
XI22698 bl<57> cbl<28> in1<72> in2<72> sl<57> vdd vss wl<72> / cell_PIM2
XI23863 bl<47> cbl<23> in1<35> in2<35> sl<47> vdd vss wl<35> / cell_PIM2
XI23862 bl<47> cbl<23> in1<36> in2<36> sl<47> vdd vss wl<36> / cell_PIM2
XI24512 bl<55> cbl<27> in1<15> in2<15> sl<55> vdd vss wl<15> / cell_PIM2
XI24511 bl<55> cbl<27> in1<16> in2<16> sl<55> vdd vss wl<16> / cell_PIM2
XI24510 bl<55> cbl<27> in1<17> in2<17> sl<55> vdd vss wl<17> / cell_PIM2
XI22688 bl<55> cbl<27> in1<72> in2<72> sl<55> vdd vss wl<72> / cell_PIM2
XI23248 bl<45> cbl<22> in1<52> in2<52> sl<45> vdd vss wl<52> / cell_PIM2
XI23247 bl<45> cbl<22> in1<51> in2<51> sl<45> vdd vss wl<51> / cell_PIM2
XI23246 bl<45> cbl<22> in1<55> in2<55> sl<45> vdd vss wl<55> / cell_PIM2
XI23245 bl<45> cbl<22> in1<54> in2<54> sl<45> vdd vss wl<54> / cell_PIM2
XI23856 bl<45> cbl<22> in1<33> in2<33> sl<45> vdd vss wl<33> / cell_PIM2
XI23855 bl<45> cbl<22> in1<32> in2<32> sl<45> vdd vss wl<32> / cell_PIM2
XI23854 bl<45> cbl<22> in1<36> in2<36> sl<45> vdd vss wl<36> / cell_PIM2
XI24504 bl<53> cbl<26> in1<14> in2<14> sl<53> vdd vss wl<14> / cell_PIM2
XI23244 bl<45> cbl<22> in1<53> in2<53> sl<45> vdd vss wl<53> / cell_PIM2
XI23853 bl<45> cbl<22> in1<35> in2<35> sl<45> vdd vss wl<35> / cell_PIM2
XI23852 bl<45> cbl<22> in1<34> in2<34> sl<45> vdd vss wl<34> / cell_PIM2
XI24502 bl<53> cbl<26> in1<17> in2<17> sl<53> vdd vss wl<17> / cell_PIM2
XI24501 bl<53> cbl<26> in1<16> in2<16> sl<53> vdd vss wl<16> / cell_PIM2
XI24500 bl<53> cbl<26> in1<15> in2<15> sl<53> vdd vss wl<15> / cell_PIM2
XI24494 bl<51> cbl<25> in1<13> in2<13> sl<51> vdd vss wl<13> / cell_PIM2
XI23846 bl<43> cbl<21> in1<32> in2<32> sl<43> vdd vss wl<32> / cell_PIM2
XI23845 bl<43> cbl<21> in1<33> in2<33> sl<43> vdd vss wl<33> / cell_PIM2
XI23844 bl<43> cbl<21> in1<34> in2<34> sl<43> vdd vss wl<34> / cell_PIM2
XI23238 bl<43> cbl<21> in1<51> in2<51> sl<43> vdd vss wl<51> / cell_PIM2
XI23237 bl<43> cbl<21> in1<52> in2<52> sl<43> vdd vss wl<52> / cell_PIM2
XI22678 bl<53> cbl<26> in1<74> in2<74> sl<53> vdd vss wl<74> / cell_PIM2
XI23236 bl<43> cbl<21> in1<53> in2<53> sl<43> vdd vss wl<53> / cell_PIM2
XI23235 bl<43> cbl<21> in1<54> in2<54> sl<43> vdd vss wl<54> / cell_PIM2
XI23234 bl<43> cbl<21> in1<55> in2<55> sl<43> vdd vss wl<55> / cell_PIM2
XI23843 bl<43> cbl<21> in1<35> in2<35> sl<43> vdd vss wl<35> / cell_PIM2
XI23842 bl<43> cbl<21> in1<36> in2<36> sl<43> vdd vss wl<36> / cell_PIM2
XI24492 bl<51> cbl<25> in1<15> in2<15> sl<51> vdd vss wl<15> / cell_PIM2
XI24491 bl<51> cbl<25> in1<16> in2<16> sl<51> vdd vss wl<16> / cell_PIM2
XI24490 bl<51> cbl<25> in1<17> in2<17> sl<51> vdd vss wl<17> / cell_PIM2
XI22668 bl<51> cbl<25> in1<72> in2<72> sl<51> vdd vss wl<72> / cell_PIM2
XI23836 bl<41> cbl<20> in1<32> in2<32> sl<41> vdd vss wl<32> / cell_PIM2
XI23835 bl<41> cbl<20> in1<33> in2<33> sl<41> vdd vss wl<33> / cell_PIM2
XI23834 bl<41> cbl<20> in1<34> in2<34> sl<41> vdd vss wl<34> / cell_PIM2
XI24484 bl<49> cbl<24> in1<14> in2<14> sl<49> vdd vss wl<14> / cell_PIM2
XI23228 bl<41> cbl<20> in1<51> in2<51> sl<41> vdd vss wl<51> / cell_PIM2
XI23227 bl<41> cbl<20> in1<52> in2<52> sl<41> vdd vss wl<52> / cell_PIM2
XI23226 bl<41> cbl<20> in1<53> in2<53> sl<41> vdd vss wl<53> / cell_PIM2
XI23225 bl<41> cbl<20> in1<54> in2<54> sl<41> vdd vss wl<54> / cell_PIM2
XI23833 bl<41> cbl<20> in1<35> in2<35> sl<41> vdd vss wl<35> / cell_PIM2
XI23832 bl<41> cbl<20> in1<36> in2<36> sl<41> vdd vss wl<36> / cell_PIM2
XI24482 bl<49> cbl<24> in1<17> in2<17> sl<49> vdd vss wl<17> / cell_PIM2
XI24481 bl<49> cbl<24> in1<16> in2<16> sl<49> vdd vss wl<16> / cell_PIM2
XI24480 bl<49> cbl<24> in1<15> in2<15> sl<49> vdd vss wl<15> / cell_PIM2
XI24474 bl<47> cbl<23> in1<13> in2<13> sl<47> vdd vss wl<13> / cell_PIM2
XI23826 bl<39> cbl<19> in1<32> in2<32> sl<39> vdd vss wl<32> / cell_PIM2
XI23825 bl<39> cbl<19> in1<33> in2<33> sl<39> vdd vss wl<33> / cell_PIM2
XI23824 bl<39> cbl<19> in1<34> in2<34> sl<39> vdd vss wl<34> / cell_PIM2
XI23224 bl<41> cbl<20> in1<55> in2<55> sl<41> vdd vss wl<55> / cell_PIM2
XI22658 bl<49> cbl<24> in1<74> in2<74> sl<49> vdd vss wl<74> / cell_PIM2
XI23218 bl<39> cbl<19> in1<51> in2<51> sl<39> vdd vss wl<51> / cell_PIM2
XI23217 bl<39> cbl<19> in1<52> in2<52> sl<39> vdd vss wl<52> / cell_PIM2
XI23823 bl<39> cbl<19> in1<35> in2<35> sl<39> vdd vss wl<35> / cell_PIM2
XI23822 bl<39> cbl<19> in1<36> in2<36> sl<39> vdd vss wl<36> / cell_PIM2
XI24472 bl<47> cbl<23> in1<15> in2<15> sl<47> vdd vss wl<15> / cell_PIM2
XI24471 bl<47> cbl<23> in1<16> in2<16> sl<47> vdd vss wl<16> / cell_PIM2
XI24470 bl<47> cbl<23> in1<17> in2<17> sl<47> vdd vss wl<17> / cell_PIM2
XI22648 bl<47> cbl<23> in1<72> in2<72> sl<47> vdd vss wl<72> / cell_PIM2
XI23216 bl<39> cbl<19> in1<53> in2<53> sl<39> vdd vss wl<53> / cell_PIM2
XI23215 bl<39> cbl<19> in1<54> in2<54> sl<39> vdd vss wl<54> / cell_PIM2
XI23214 bl<39> cbl<19> in1<55> in2<55> sl<39> vdd vss wl<55> / cell_PIM2
XI23816 bl<37> cbl<18> in1<33> in2<33> sl<37> vdd vss wl<33> / cell_PIM2
XI23815 bl<37> cbl<18> in1<32> in2<32> sl<37> vdd vss wl<32> / cell_PIM2
XI23814 bl<37> cbl<18> in1<36> in2<36> sl<37> vdd vss wl<36> / cell_PIM2
XI24464 bl<45> cbl<22> in1<14> in2<14> sl<45> vdd vss wl<14> / cell_PIM2
XI23813 bl<37> cbl<18> in1<35> in2<35> sl<37> vdd vss wl<35> / cell_PIM2
XI23812 bl<37> cbl<18> in1<34> in2<34> sl<37> vdd vss wl<34> / cell_PIM2
XI24462 bl<45> cbl<22> in1<17> in2<17> sl<45> vdd vss wl<17> / cell_PIM2
XI24461 bl<45> cbl<22> in1<16> in2<16> sl<45> vdd vss wl<16> / cell_PIM2
XI24460 bl<45> cbl<22> in1<15> in2<15> sl<45> vdd vss wl<15> / cell_PIM2
XI24454 bl<43> cbl<21> in1<13> in2<13> sl<43> vdd vss wl<13> / cell_PIM2
XI23806 bl<35> cbl<17> in1<32> in2<32> sl<35> vdd vss wl<32> / cell_PIM2
XI23805 bl<35> cbl<17> in1<33> in2<33> sl<35> vdd vss wl<33> / cell_PIM2
XI23804 bl<35> cbl<17> in1<34> in2<34> sl<35> vdd vss wl<34> / cell_PIM2
XI23208 bl<37> cbl<18> in1<52> in2<52> sl<37> vdd vss wl<52> / cell_PIM2
XI23207 bl<37> cbl<18> in1<51> in2<51> sl<37> vdd vss wl<51> / cell_PIM2
XI23206 bl<37> cbl<18> in1<55> in2<55> sl<37> vdd vss wl<55> / cell_PIM2
XI23205 bl<37> cbl<18> in1<54> in2<54> sl<37> vdd vss wl<54> / cell_PIM2
XI22638 bl<45> cbl<22> in1<74> in2<74> sl<45> vdd vss wl<74> / cell_PIM2
XI23204 bl<37> cbl<18> in1<53> in2<53> sl<37> vdd vss wl<53> / cell_PIM2
XI23803 bl<35> cbl<17> in1<35> in2<35> sl<35> vdd vss wl<35> / cell_PIM2
XI23802 bl<35> cbl<17> in1<36> in2<36> sl<35> vdd vss wl<36> / cell_PIM2
XI24452 bl<43> cbl<21> in1<15> in2<15> sl<43> vdd vss wl<15> / cell_PIM2
XI24451 bl<43> cbl<21> in1<16> in2<16> sl<43> vdd vss wl<16> / cell_PIM2
XI24450 bl<43> cbl<21> in1<17> in2<17> sl<43> vdd vss wl<17> / cell_PIM2
XI22628 bl<43> cbl<21> in1<72> in2<72> sl<43> vdd vss wl<72> / cell_PIM2
XI23198 bl<35> cbl<17> in1<51> in2<51> sl<35> vdd vss wl<51> / cell_PIM2
XI23197 bl<35> cbl<17> in1<52> in2<52> sl<35> vdd vss wl<52> / cell_PIM2
XI23796 bl<33> cbl<16> in1<33> in2<33> sl<33> vdd vss wl<33> / cell_PIM2
XI23795 bl<33> cbl<16> in1<32> in2<32> sl<33> vdd vss wl<32> / cell_PIM2
XI23794 bl<33> cbl<16> in1<36> in2<36> sl<33> vdd vss wl<36> / cell_PIM2
XI24444 bl<41> cbl<20> in1<13> in2<13> sl<41> vdd vss wl<13> / cell_PIM2
XI23196 bl<35> cbl<17> in1<53> in2<53> sl<35> vdd vss wl<53> / cell_PIM2
XI23195 bl<35> cbl<17> in1<54> in2<54> sl<35> vdd vss wl<54> / cell_PIM2
XI23194 bl<35> cbl<17> in1<55> in2<55> sl<35> vdd vss wl<55> / cell_PIM2
XI23793 bl<33> cbl<16> in1<35> in2<35> sl<33> vdd vss wl<35> / cell_PIM2
XI23792 bl<33> cbl<16> in1<34> in2<34> sl<33> vdd vss wl<34> / cell_PIM2
XI24442 bl<41> cbl<20> in1<15> in2<15> sl<41> vdd vss wl<15> / cell_PIM2
XI24441 bl<41> cbl<20> in1<16> in2<16> sl<41> vdd vss wl<16> / cell_PIM2
XI24440 bl<41> cbl<20> in1<17> in2<17> sl<41> vdd vss wl<17> / cell_PIM2
XI24434 bl<39> cbl<19> in1<13> in2<13> sl<39> vdd vss wl<13> / cell_PIM2
XI23786 bl<63> cbl<31> in1<37> in2<37> sl<63> vdd vss wl<37> / cell_PIM2
XI23785 bl<63> cbl<31> in1<38> in2<38> sl<63> vdd vss wl<38> / cell_PIM2
XI23784 bl<63> cbl<31> in1<39> in2<39> sl<63> vdd vss wl<39> / cell_PIM2
XI22618 bl<41> cbl<20> in1<72> in2<72> sl<41> vdd vss wl<72> / cell_PIM2
XI23188 bl<33> cbl<16> in1<52> in2<52> sl<33> vdd vss wl<52> / cell_PIM2
XI23187 bl<33> cbl<16> in1<51> in2<51> sl<33> vdd vss wl<51> / cell_PIM2
XI23186 bl<33> cbl<16> in1<55> in2<55> sl<33> vdd vss wl<55> / cell_PIM2
XI23185 bl<33> cbl<16> in1<54> in2<54> sl<33> vdd vss wl<54> / cell_PIM2
XI23783 bl<63> cbl<31> in1<40> in2<40> sl<63> vdd vss wl<40> / cell_PIM2
XI24432 bl<39> cbl<19> in1<15> in2<15> sl<39> vdd vss wl<15> / cell_PIM2
XI24431 bl<39> cbl<19> in1<16> in2<16> sl<39> vdd vss wl<16> / cell_PIM2
XI24430 bl<39> cbl<19> in1<17> in2<17> sl<39> vdd vss wl<17> / cell_PIM2
XI22608 bl<39> cbl<19> in1<72> in2<72> sl<39> vdd vss wl<72> / cell_PIM2
XI23184 bl<33> cbl<16> in1<53> in2<53> sl<33> vdd vss wl<53> / cell_PIM2
XI23778 bl<61> cbl<30> in1<38> in2<38> sl<61> vdd vss wl<38> / cell_PIM2
XI23777 bl<61> cbl<30> in1<37> in2<37> sl<61> vdd vss wl<37> / cell_PIM2
XI23776 bl<61> cbl<30> in1<40> in2<40> sl<61> vdd vss wl<40> / cell_PIM2
XI23775 bl<61> cbl<30> in1<39> in2<39> sl<61> vdd vss wl<39> / cell_PIM2
XI24424 bl<37> cbl<18> in1<14> in2<14> sl<37> vdd vss wl<14> / cell_PIM2
XI23178 bl<63> cbl<31> in1<56> in2<56> sl<63> vdd vss wl<56> / cell_PIM2
XI23177 bl<63> cbl<31> in1<57> in2<57> sl<63> vdd vss wl<57> / cell_PIM2
XI23770 bl<59> cbl<29> in1<37> in2<37> sl<59> vdd vss wl<37> / cell_PIM2
XI23769 bl<59> cbl<29> in1<38> in2<38> sl<59> vdd vss wl<38> / cell_PIM2
XI24422 bl<37> cbl<18> in1<17> in2<17> sl<37> vdd vss wl<17> / cell_PIM2
XI24421 bl<37> cbl<18> in1<16> in2<16> sl<37> vdd vss wl<16> / cell_PIM2
XI24420 bl<37> cbl<18> in1<15> in2<15> sl<37> vdd vss wl<15> / cell_PIM2
XI24414 bl<35> cbl<17> in1<13> in2<13> sl<35> vdd vss wl<13> / cell_PIM2
XI23768 bl<59> cbl<29> in1<39> in2<39> sl<59> vdd vss wl<39> / cell_PIM2
XI23767 bl<59> cbl<29> in1<40> in2<40> sl<59> vdd vss wl<40> / cell_PIM2
XI23176 bl<63> cbl<31> in1<58> in2<58> sl<63> vdd vss wl<58> / cell_PIM2
XI23175 bl<63> cbl<31> in1<59> in2<59> sl<63> vdd vss wl<59> / cell_PIM2
XI23174 bl<63> cbl<31> in1<60> in2<60> sl<63> vdd vss wl<60> / cell_PIM2
XI22598 bl<37> cbl<18> in1<74> in2<74> sl<37> vdd vss wl<74> / cell_PIM2
XI23762 bl<57> cbl<28> in1<37> in2<37> sl<57> vdd vss wl<37> / cell_PIM2
XI23761 bl<57> cbl<28> in1<38> in2<38> sl<57> vdd vss wl<38> / cell_PIM2
XI23760 bl<57> cbl<28> in1<39> in2<39> sl<57> vdd vss wl<39> / cell_PIM2
XI23759 bl<57> cbl<28> in1<40> in2<40> sl<57> vdd vss wl<40> / cell_PIM2
XI24412 bl<35> cbl<17> in1<15> in2<15> sl<35> vdd vss wl<15> / cell_PIM2
XI24411 bl<35> cbl<17> in1<16> in2<16> sl<35> vdd vss wl<16> / cell_PIM2
XI24410 bl<35> cbl<17> in1<17> in2<17> sl<35> vdd vss wl<17> / cell_PIM2
XI22588 bl<35> cbl<17> in1<72> in2<72> sl<35> vdd vss wl<72> / cell_PIM2
XI23168 bl<61> cbl<30> in1<57> in2<57> sl<61> vdd vss wl<57> / cell_PIM2
XI23167 bl<61> cbl<30> in1<56> in2<56> sl<61> vdd vss wl<56> / cell_PIM2
XI23166 bl<61> cbl<30> in1<60> in2<60> sl<61> vdd vss wl<60> / cell_PIM2
XI23165 bl<61> cbl<30> in1<59> in2<59> sl<61> vdd vss wl<59> / cell_PIM2
XI23754 bl<55> cbl<27> in1<37> in2<37> sl<55> vdd vss wl<37> / cell_PIM2
XI24404 bl<33> cbl<16> in1<14> in2<14> sl<33> vdd vss wl<14> / cell_PIM2
XI23164 bl<61> cbl<30> in1<58> in2<58> sl<61> vdd vss wl<58> / cell_PIM2
XI23753 bl<55> cbl<27> in1<38> in2<38> sl<55> vdd vss wl<38> / cell_PIM2
XI23752 bl<55> cbl<27> in1<39> in2<39> sl<55> vdd vss wl<39> / cell_PIM2
XI23751 bl<55> cbl<27> in1<40> in2<40> sl<55> vdd vss wl<40> / cell_PIM2
XI24402 bl<33> cbl<16> in1<17> in2<17> sl<33> vdd vss wl<17> / cell_PIM2
XI24401 bl<33> cbl<16> in1<16> in2<16> sl<33> vdd vss wl<16> / cell_PIM2
XI24400 bl<33> cbl<16> in1<15> in2<15> sl<33> vdd vss wl<15> / cell_PIM2
XI24394 bl<63> cbl<31> in1<18> in2<18> sl<63> vdd vss wl<18> / cell_PIM2
XI23746 bl<53> cbl<26> in1<38> in2<38> sl<53> vdd vss wl<38> / cell_PIM2
XI23745 bl<53> cbl<26> in1<37> in2<37> sl<53> vdd vss wl<37> / cell_PIM2
XI23744 bl<53> cbl<26> in1<40> in2<40> sl<53> vdd vss wl<40> / cell_PIM2
XI23158 bl<59> cbl<29> in1<56> in2<56> sl<59> vdd vss wl<56> / cell_PIM2
XI23157 bl<59> cbl<29> in1<57> in2<57> sl<59> vdd vss wl<57> / cell_PIM2
XI22578 bl<33> cbl<16> in1<74> in2<74> sl<33> vdd vss wl<74> / cell_PIM2
XI23156 bl<59> cbl<29> in1<58> in2<58> sl<59> vdd vss wl<58> / cell_PIM2
XI23155 bl<59> cbl<29> in1<59> in2<59> sl<59> vdd vss wl<59> / cell_PIM2
XI23154 bl<59> cbl<29> in1<60> in2<60> sl<59> vdd vss wl<60> / cell_PIM2
XI23743 bl<53> cbl<26> in1<39> in2<39> sl<53> vdd vss wl<39> / cell_PIM2
XI24392 bl<63> cbl<31> in1<20> in2<20> sl<63> vdd vss wl<20> / cell_PIM2
XI24391 bl<63> cbl<31> in1<21> in2<21> sl<63> vdd vss wl<21> / cell_PIM2
XI22568 bl<63> cbl<31> in1<77> in2<77> sl<63> vdd vss wl<77> / cell_PIM2
XI23738 bl<51> cbl<25> in1<37> in2<37> sl<51> vdd vss wl<37> / cell_PIM2
XI23737 bl<51> cbl<25> in1<38> in2<38> sl<51> vdd vss wl<38> / cell_PIM2
XI23736 bl<51> cbl<25> in1<39> in2<39> sl<51> vdd vss wl<39> / cell_PIM2
XI23735 bl<51> cbl<25> in1<40> in2<40> sl<51> vdd vss wl<40> / cell_PIM2
XI24386 bl<61> cbl<30> in1<19> in2<19> sl<61> vdd vss wl<19> / cell_PIM2
XI24385 bl<61> cbl<30> in1<18> in2<18> sl<61> vdd vss wl<18> / cell_PIM2
XI24384 bl<61> cbl<30> in1<21> in2<21> sl<61> vdd vss wl<21> / cell_PIM2
XI21583 bl<49> cbl<24> in1<106> in2<106> sl<49> vdd vss wl<106> / cell_PIM2
XI22232 bl<53> cbl<26> in1<86> in2<86> sl<53> vdd vss wl<86> / cell_PIM2
XI22231 bl<53> cbl<26> in1<85> in2<85> sl<53> vdd vss wl<85> / cell_PIM2
XI22230 bl<53> cbl<26> in1<84> in2<84> sl<53> vdd vss wl<84> / cell_PIM2
XI22229 bl<53> cbl<26> in1<88> in2<88> sl<53> vdd vss wl<88> / cell_PIM2
XI22880 bl<61> cbl<30> in1<67> in2<67> sl<61> vdd vss wl<67> / cell_PIM2
XI22879 bl<61> cbl<30> in1<66> in2<66> sl<61> vdd vss wl<66> / cell_PIM2
XI22877 bl<61> cbl<30> in1<69> in2<69> sl<61> vdd vss wl<69> / cell_PIM2
XI22876 bl<61> cbl<30> in1<68> in2<68> sl<61> vdd vss wl<68> / cell_PIM2
XI22228 bl<53> cbl<26> in1<87> in2<87> sl<53> vdd vss wl<87> / cell_PIM2
XI21578 bl<47> cbl<23> in1<104> in2<104> sl<47> vdd vss wl<104> / cell_PIM2
XI21577 bl<47> cbl<23> in1<105> in2<105> sl<47> vdd vss wl<105> / cell_PIM2
XI21576 bl<47> cbl<23> in1<106> in2<106> sl<47> vdd vss wl<106> / cell_PIM2
XI21575 bl<47> cbl<23> in1<107> in2<107> sl<47> vdd vss wl<107> / cell_PIM2
XI21570 bl<45> cbl<22> in1<105> in2<105> sl<45> vdd vss wl<105> / cell_PIM2
XI21569 bl<45> cbl<22> in1<104> in2<104> sl<45> vdd vss wl<104> / cell_PIM2
XI22222 bl<51> cbl<25> in1<84> in2<84> sl<51> vdd vss wl<84> / cell_PIM2
XI22221 bl<51> cbl<25> in1<85> in2<85> sl<51> vdd vss wl<85> / cell_PIM2
XI22220 bl<51> cbl<25> in1<86> in2<86> sl<51> vdd vss wl<86> / cell_PIM2
XI22219 bl<51> cbl<25> in1<87> in2<87> sl<51> vdd vss wl<87> / cell_PIM2
XI22870 bl<59> cbl<29> in1<65> in2<65> sl<59> vdd vss wl<65> / cell_PIM2
XI22869 bl<59> cbl<29> in1<66> in2<66> sl<59> vdd vss wl<66> / cell_PIM2
XI21568 bl<45> cbl<22> in1<107> in2<107> sl<45> vdd vss wl<107> / cell_PIM2
XI21567 bl<45> cbl<22> in1<106> in2<106> sl<45> vdd vss wl<106> / cell_PIM2
XI22218 bl<51> cbl<25> in1<88> in2<88> sl<51> vdd vss wl<88> / cell_PIM2
XI22867 bl<59> cbl<29> in1<68> in2<68> sl<59> vdd vss wl<68> / cell_PIM2
XI22866 bl<59> cbl<29> in1<69> in2<69> sl<59> vdd vss wl<69> / cell_PIM2
XI21562 bl<43> cbl<21> in1<104> in2<104> sl<43> vdd vss wl<104> / cell_PIM2
XI21561 bl<43> cbl<21> in1<105> in2<105> sl<43> vdd vss wl<105> / cell_PIM2
XI21560 bl<43> cbl<21> in1<106> in2<106> sl<43> vdd vss wl<106> / cell_PIM2
XI21559 bl<43> cbl<21> in1<107> in2<107> sl<43> vdd vss wl<107> / cell_PIM2
XI22212 bl<49> cbl<24> in1<86> in2<86> sl<49> vdd vss wl<86> / cell_PIM2
XI22211 bl<49> cbl<24> in1<85> in2<85> sl<49> vdd vss wl<85> / cell_PIM2
XI22210 bl<49> cbl<24> in1<84> in2<84> sl<49> vdd vss wl<84> / cell_PIM2
XI22209 bl<49> cbl<24> in1<88> in2<88> sl<49> vdd vss wl<88> / cell_PIM2
XI22860 bl<57> cbl<28> in1<65> in2<65> sl<57> vdd vss wl<65> / cell_PIM2
XI22859 bl<57> cbl<28> in1<66> in2<66> sl<57> vdd vss wl<66> / cell_PIM2
XI22857 bl<57> cbl<28> in1<68> in2<68> sl<57> vdd vss wl<68> / cell_PIM2
XI22856 bl<57> cbl<28> in1<69> in2<69> sl<57> vdd vss wl<69> / cell_PIM2
XI22208 bl<49> cbl<24> in1<87> in2<87> sl<49> vdd vss wl<87> / cell_PIM2
XI21554 bl<41> cbl<20> in1<104> in2<104> sl<41> vdd vss wl<104> / cell_PIM2
XI21553 bl<41> cbl<20> in1<105> in2<105> sl<41> vdd vss wl<105> / cell_PIM2
XI21552 bl<41> cbl<20> in1<106> in2<106> sl<41> vdd vss wl<106> / cell_PIM2
XI21551 bl<41> cbl<20> in1<107> in2<107> sl<41> vdd vss wl<107> / cell_PIM2
XI22202 bl<47> cbl<23> in1<84> in2<84> sl<47> vdd vss wl<84> / cell_PIM2
XI22201 bl<47> cbl<23> in1<85> in2<85> sl<47> vdd vss wl<85> / cell_PIM2
XI22200 bl<47> cbl<23> in1<86> in2<86> sl<47> vdd vss wl<86> / cell_PIM2
XI22199 bl<47> cbl<23> in1<87> in2<87> sl<47> vdd vss wl<87> / cell_PIM2
XI22850 bl<55> cbl<27> in1<65> in2<65> sl<55> vdd vss wl<65> / cell_PIM2
XI22849 bl<55> cbl<27> in1<66> in2<66> sl<55> vdd vss wl<66> / cell_PIM2
XI21546 bl<39> cbl<19> in1<104> in2<104> sl<39> vdd vss wl<104> / cell_PIM2
XI21545 bl<39> cbl<19> in1<105> in2<105> sl<39> vdd vss wl<105> / cell_PIM2
XI21544 bl<39> cbl<19> in1<106> in2<106> sl<39> vdd vss wl<106> / cell_PIM2
XI22198 bl<47> cbl<23> in1<88> in2<88> sl<47> vdd vss wl<88> / cell_PIM2
XI22847 bl<55> cbl<27> in1<68> in2<68> sl<55> vdd vss wl<68> / cell_PIM2
XI22846 bl<55> cbl<27> in1<69> in2<69> sl<55> vdd vss wl<69> / cell_PIM2
XI21543 bl<39> cbl<19> in1<107> in2<107> sl<39> vdd vss wl<107> / cell_PIM2
XI22192 bl<45> cbl<22> in1<86> in2<86> sl<45> vdd vss wl<86> / cell_PIM2
XI22191 bl<45> cbl<22> in1<85> in2<85> sl<45> vdd vss wl<85> / cell_PIM2
XI22190 bl<45> cbl<22> in1<84> in2<84> sl<45> vdd vss wl<84> / cell_PIM2
XI22189 bl<45> cbl<22> in1<88> in2<88> sl<45> vdd vss wl<88> / cell_PIM2
XI22840 bl<53> cbl<26> in1<67> in2<67> sl<53> vdd vss wl<67> / cell_PIM2
XI22839 bl<53> cbl<26> in1<66> in2<66> sl<53> vdd vss wl<66> / cell_PIM2
XI22837 bl<53> cbl<26> in1<69> in2<69> sl<53> vdd vss wl<69> / cell_PIM2
XI22836 bl<53> cbl<26> in1<68> in2<68> sl<53> vdd vss wl<68> / cell_PIM2
XI22188 bl<45> cbl<22> in1<87> in2<87> sl<45> vdd vss wl<87> / cell_PIM2
XI21538 bl<37> cbl<18> in1<105> in2<105> sl<37> vdd vss wl<105> / cell_PIM2
XI21537 bl<37> cbl<18> in1<104> in2<104> sl<37> vdd vss wl<104> / cell_PIM2
XI21536 bl<37> cbl<18> in1<107> in2<107> sl<37> vdd vss wl<107> / cell_PIM2
XI21535 bl<37> cbl<18> in1<106> in2<106> sl<37> vdd vss wl<106> / cell_PIM2
XI21530 bl<35> cbl<17> in1<104> in2<104> sl<35> vdd vss wl<104> / cell_PIM2
XI21529 bl<35> cbl<17> in1<105> in2<105> sl<35> vdd vss wl<105> / cell_PIM2
XI22182 bl<43> cbl<21> in1<84> in2<84> sl<43> vdd vss wl<84> / cell_PIM2
XI22181 bl<43> cbl<21> in1<85> in2<85> sl<43> vdd vss wl<85> / cell_PIM2
XI22180 bl<43> cbl<21> in1<86> in2<86> sl<43> vdd vss wl<86> / cell_PIM2
XI22179 bl<43> cbl<21> in1<87> in2<87> sl<43> vdd vss wl<87> / cell_PIM2
XI22830 bl<51> cbl<25> in1<65> in2<65> sl<51> vdd vss wl<65> / cell_PIM2
XI22829 bl<51> cbl<25> in1<66> in2<66> sl<51> vdd vss wl<66> / cell_PIM2
XI21528 bl<35> cbl<17> in1<106> in2<106> sl<35> vdd vss wl<106> / cell_PIM2
XI21527 bl<35> cbl<17> in1<107> in2<107> sl<35> vdd vss wl<107> / cell_PIM2
XI22178 bl<43> cbl<21> in1<88> in2<88> sl<43> vdd vss wl<88> / cell_PIM2
XI22827 bl<51> cbl<25> in1<68> in2<68> sl<51> vdd vss wl<68> / cell_PIM2
XI22826 bl<51> cbl<25> in1<69> in2<69> sl<51> vdd vss wl<69> / cell_PIM2
XI21522 bl<33> cbl<16> in1<105> in2<105> sl<33> vdd vss wl<105> / cell_PIM2
XI21521 bl<33> cbl<16> in1<104> in2<104> sl<33> vdd vss wl<104> / cell_PIM2
XI21520 bl<33> cbl<16> in1<107> in2<107> sl<33> vdd vss wl<107> / cell_PIM2
XI21519 bl<33> cbl<16> in1<106> in2<106> sl<33> vdd vss wl<106> / cell_PIM2
XI22172 bl<41> cbl<20> in1<84> in2<84> sl<41> vdd vss wl<84> / cell_PIM2
XI22171 bl<41> cbl<20> in1<85> in2<85> sl<41> vdd vss wl<85> / cell_PIM2
XI22170 bl<41> cbl<20> in1<86> in2<86> sl<41> vdd vss wl<86> / cell_PIM2
XI22169 bl<41> cbl<20> in1<87> in2<87> sl<41> vdd vss wl<87> / cell_PIM2
XI22820 bl<49> cbl<24> in1<67> in2<67> sl<49> vdd vss wl<67> / cell_PIM2
XI22819 bl<49> cbl<24> in1<66> in2<66> sl<49> vdd vss wl<66> / cell_PIM2
XI22817 bl<49> cbl<24> in1<69> in2<69> sl<49> vdd vss wl<69> / cell_PIM2
XI22816 bl<49> cbl<24> in1<68> in2<68> sl<49> vdd vss wl<68> / cell_PIM2
XI22168 bl<41> cbl<20> in1<88> in2<88> sl<41> vdd vss wl<88> / cell_PIM2
XI21514 bl<63> cbl<31> in1<108> in2<108> sl<63> vdd vss wl<108> / cell_PIM2
XI21513 bl<63> cbl<31> in1<109> in2<109> sl<63> vdd vss wl<109> / cell_PIM2
XI21512 bl<63> cbl<31> in1<110> in2<110> sl<63> vdd vss wl<110> / cell_PIM2
XI21511 bl<63> cbl<31> in1<111> in2<111> sl<63> vdd vss wl<111> / cell_PIM2
XI21510 bl<63> cbl<31> in1<112> in2<112> sl<63> vdd vss wl<112> / cell_PIM2
XI22162 bl<39> cbl<19> in1<84> in2<84> sl<39> vdd vss wl<84> / cell_PIM2
XI22161 bl<39> cbl<19> in1<85> in2<85> sl<39> vdd vss wl<85> / cell_PIM2
XI22160 bl<39> cbl<19> in1<86> in2<86> sl<39> vdd vss wl<86> / cell_PIM2
XI22159 bl<39> cbl<19> in1<87> in2<87> sl<39> vdd vss wl<87> / cell_PIM2
XI22810 bl<47> cbl<23> in1<65> in2<65> sl<47> vdd vss wl<65> / cell_PIM2
XI22809 bl<47> cbl<23> in1<66> in2<66> sl<47> vdd vss wl<66> / cell_PIM2
XI21504 bl<61> cbl<30> in1<110> in2<110> sl<61> vdd vss wl<110> / cell_PIM2
XI22158 bl<39> cbl<19> in1<88> in2<88> sl<39> vdd vss wl<88> / cell_PIM2
XI22807 bl<47> cbl<23> in1<68> in2<68> sl<47> vdd vss wl<68> / cell_PIM2
XI22806 bl<47> cbl<23> in1<69> in2<69> sl<47> vdd vss wl<69> / cell_PIM2
XI21503 bl<61> cbl<30> in1<109> in2<109> sl<61> vdd vss wl<109> / cell_PIM2
XI21502 bl<61> cbl<30> in1<108> in2<108> sl<61> vdd vss wl<108> / cell_PIM2
XI21501 bl<61> cbl<30> in1<112> in2<112> sl<61> vdd vss wl<112> / cell_PIM2
XI21500 bl<61> cbl<30> in1<111> in2<111> sl<61> vdd vss wl<111> / cell_PIM2
XI22152 bl<37> cbl<18> in1<86> in2<86> sl<37> vdd vss wl<86> / cell_PIM2
XI22151 bl<37> cbl<18> in1<85> in2<85> sl<37> vdd vss wl<85> / cell_PIM2
XI22150 bl<37> cbl<18> in1<84> in2<84> sl<37> vdd vss wl<84> / cell_PIM2
XI22149 bl<37> cbl<18> in1<88> in2<88> sl<37> vdd vss wl<88> / cell_PIM2
XI22800 bl<45> cbl<22> in1<67> in2<67> sl<45> vdd vss wl<67> / cell_PIM2
XI22799 bl<45> cbl<22> in1<66> in2<66> sl<45> vdd vss wl<66> / cell_PIM2
XI22797 bl<45> cbl<22> in1<69> in2<69> sl<45> vdd vss wl<69> / cell_PIM2
XI22796 bl<45> cbl<22> in1<68> in2<68> sl<45> vdd vss wl<68> / cell_PIM2
XI22148 bl<37> cbl<18> in1<87> in2<87> sl<37> vdd vss wl<87> / cell_PIM2
XI21494 bl<59> cbl<29> in1<108> in2<108> sl<59> vdd vss wl<108> / cell_PIM2
XI21493 bl<59> cbl<29> in1<109> in2<109> sl<59> vdd vss wl<109> / cell_PIM2
XI21492 bl<59> cbl<29> in1<110> in2<110> sl<59> vdd vss wl<110> / cell_PIM2
XI21491 bl<59> cbl<29> in1<111> in2<111> sl<59> vdd vss wl<111> / cell_PIM2
XI21490 bl<59> cbl<29> in1<112> in2<112> sl<59> vdd vss wl<112> / cell_PIM2
XI22142 bl<35> cbl<17> in1<84> in2<84> sl<35> vdd vss wl<84> / cell_PIM2
XI22141 bl<35> cbl<17> in1<85> in2<85> sl<35> vdd vss wl<85> / cell_PIM2
XI22140 bl<35> cbl<17> in1<86> in2<86> sl<35> vdd vss wl<86> / cell_PIM2
XI22139 bl<35> cbl<17> in1<87> in2<87> sl<35> vdd vss wl<87> / cell_PIM2
XI22790 bl<43> cbl<21> in1<65> in2<65> sl<43> vdd vss wl<65> / cell_PIM2
XI22789 bl<43> cbl<21> in1<66> in2<66> sl<43> vdd vss wl<66> / cell_PIM2
XI21484 bl<57> cbl<28> in1<108> in2<108> sl<57> vdd vss wl<108> / cell_PIM2
XI22138 bl<35> cbl<17> in1<88> in2<88> sl<35> vdd vss wl<88> / cell_PIM2
XI22787 bl<43> cbl<21> in1<68> in2<68> sl<43> vdd vss wl<68> / cell_PIM2
XI22786 bl<43> cbl<21> in1<69> in2<69> sl<43> vdd vss wl<69> / cell_PIM2
XI21483 bl<57> cbl<28> in1<109> in2<109> sl<57> vdd vss wl<109> / cell_PIM2
XI21482 bl<57> cbl<28> in1<110> in2<110> sl<57> vdd vss wl<110> / cell_PIM2
XI21481 bl<57> cbl<28> in1<111> in2<111> sl<57> vdd vss wl<111> / cell_PIM2
XI21480 bl<57> cbl<28> in1<112> in2<112> sl<57> vdd vss wl<112> / cell_PIM2
XI22132 bl<33> cbl<16> in1<86> in2<86> sl<33> vdd vss wl<86> / cell_PIM2
XI22131 bl<33> cbl<16> in1<85> in2<85> sl<33> vdd vss wl<85> / cell_PIM2
XI22130 bl<33> cbl<16> in1<84> in2<84> sl<33> vdd vss wl<84> / cell_PIM2
XI22129 bl<33> cbl<16> in1<88> in2<88> sl<33> vdd vss wl<88> / cell_PIM2
XI22780 bl<41> cbl<20> in1<65> in2<65> sl<41> vdd vss wl<65> / cell_PIM2
XI22779 bl<41> cbl<20> in1<66> in2<66> sl<41> vdd vss wl<66> / cell_PIM2
XI22777 bl<41> cbl<20> in1<68> in2<68> sl<41> vdd vss wl<68> / cell_PIM2
XI22776 bl<41> cbl<20> in1<69> in2<69> sl<41> vdd vss wl<69> / cell_PIM2
XI22128 bl<33> cbl<16> in1<87> in2<87> sl<33> vdd vss wl<87> / cell_PIM2
XI21474 bl<55> cbl<27> in1<108> in2<108> sl<55> vdd vss wl<108> / cell_PIM2
XI21473 bl<55> cbl<27> in1<109> in2<109> sl<55> vdd vss wl<109> / cell_PIM2
XI21472 bl<55> cbl<27> in1<110> in2<110> sl<55> vdd vss wl<110> / cell_PIM2
XI21471 bl<55> cbl<27> in1<111> in2<111> sl<55> vdd vss wl<111> / cell_PIM2
XI21470 bl<55> cbl<27> in1<112> in2<112> sl<55> vdd vss wl<112> / cell_PIM2
XI22122 bl<63> cbl<31> in1<89> in2<89> sl<63> vdd vss wl<89> / cell_PIM2
XI22121 bl<63> cbl<31> in1<90> in2<90> sl<63> vdd vss wl<90> / cell_PIM2
XI22120 bl<63> cbl<31> in1<91> in2<91> sl<63> vdd vss wl<91> / cell_PIM2
XI22119 bl<63> cbl<31> in1<92> in2<92> sl<63> vdd vss wl<92> / cell_PIM2
XI22770 bl<39> cbl<19> in1<65> in2<65> sl<39> vdd vss wl<65> / cell_PIM2
XI22769 bl<39> cbl<19> in1<66> in2<66> sl<39> vdd vss wl<66> / cell_PIM2
XI21464 bl<53> cbl<26> in1<110> in2<110> sl<53> vdd vss wl<110> / cell_PIM2
XI22118 bl<63> cbl<31> in1<93> in2<93> sl<63> vdd vss wl<93> / cell_PIM2
XI22767 bl<39> cbl<19> in1<68> in2<68> sl<39> vdd vss wl<68> / cell_PIM2
XI22766 bl<39> cbl<19> in1<69> in2<69> sl<39> vdd vss wl<69> / cell_PIM2
XI21463 bl<53> cbl<26> in1<109> in2<109> sl<53> vdd vss wl<109> / cell_PIM2
XI21462 bl<53> cbl<26> in1<108> in2<108> sl<53> vdd vss wl<108> / cell_PIM2
XI21461 bl<53> cbl<26> in1<112> in2<112> sl<53> vdd vss wl<112> / cell_PIM2
XI21460 bl<53> cbl<26> in1<111> in2<111> sl<53> vdd vss wl<111> / cell_PIM2
XI22112 bl<61> cbl<30> in1<91> in2<91> sl<61> vdd vss wl<91> / cell_PIM2
XI22111 bl<61> cbl<30> in1<90> in2<90> sl<61> vdd vss wl<90> / cell_PIM2
XI22110 bl<61> cbl<30> in1<89> in2<89> sl<61> vdd vss wl<89> / cell_PIM2
XI22109 bl<61> cbl<30> in1<93> in2<93> sl<61> vdd vss wl<93> / cell_PIM2
XI22760 bl<37> cbl<18> in1<67> in2<67> sl<37> vdd vss wl<67> / cell_PIM2
XI22759 bl<37> cbl<18> in1<66> in2<66> sl<37> vdd vss wl<66> / cell_PIM2
XI22757 bl<37> cbl<18> in1<69> in2<69> sl<37> vdd vss wl<69> / cell_PIM2
XI22756 bl<37> cbl<18> in1<68> in2<68> sl<37> vdd vss wl<68> / cell_PIM2
XI22108 bl<61> cbl<30> in1<92> in2<92> sl<61> vdd vss wl<92> / cell_PIM2
XI21454 bl<51> cbl<25> in1<108> in2<108> sl<51> vdd vss wl<108> / cell_PIM2
XI21453 bl<51> cbl<25> in1<109> in2<109> sl<51> vdd vss wl<109> / cell_PIM2
XI21452 bl<51> cbl<25> in1<110> in2<110> sl<51> vdd vss wl<110> / cell_PIM2
XI21451 bl<51> cbl<25> in1<111> in2<111> sl<51> vdd vss wl<111> / cell_PIM2
XI21450 bl<51> cbl<25> in1<112> in2<112> sl<51> vdd vss wl<112> / cell_PIM2
XI22102 bl<59> cbl<29> in1<89> in2<89> sl<59> vdd vss wl<89> / cell_PIM2
XI22101 bl<59> cbl<29> in1<90> in2<90> sl<59> vdd vss wl<90> / cell_PIM2
XI22100 bl<59> cbl<29> in1<91> in2<91> sl<59> vdd vss wl<91> / cell_PIM2
XI22099 bl<59> cbl<29> in1<92> in2<92> sl<59> vdd vss wl<92> / cell_PIM2
XI22750 bl<35> cbl<17> in1<65> in2<65> sl<35> vdd vss wl<65> / cell_PIM2
XI22749 bl<35> cbl<17> in1<66> in2<66> sl<35> vdd vss wl<66> / cell_PIM2
XI21444 bl<49> cbl<24> in1<110> in2<110> sl<49> vdd vss wl<110> / cell_PIM2
XI22098 bl<59> cbl<29> in1<93> in2<93> sl<59> vdd vss wl<93> / cell_PIM2
XI22747 bl<35> cbl<17> in1<68> in2<68> sl<35> vdd vss wl<68> / cell_PIM2
XI22746 bl<35> cbl<17> in1<69> in2<69> sl<35> vdd vss wl<69> / cell_PIM2
XI21443 bl<49> cbl<24> in1<109> in2<109> sl<49> vdd vss wl<109> / cell_PIM2
XI21442 bl<49> cbl<24> in1<108> in2<108> sl<49> vdd vss wl<108> / cell_PIM2
XI21441 bl<49> cbl<24> in1<112> in2<112> sl<49> vdd vss wl<112> / cell_PIM2
XI21440 bl<49> cbl<24> in1<111> in2<111> sl<49> vdd vss wl<111> / cell_PIM2
XI22092 bl<57> cbl<28> in1<89> in2<89> sl<57> vdd vss wl<89> / cell_PIM2
XI22091 bl<57> cbl<28> in1<90> in2<90> sl<57> vdd vss wl<90> / cell_PIM2
XI22090 bl<57> cbl<28> in1<91> in2<91> sl<57> vdd vss wl<91> / cell_PIM2
XI22089 bl<57> cbl<28> in1<92> in2<92> sl<57> vdd vss wl<92> / cell_PIM2
XI22740 bl<33> cbl<16> in1<67> in2<67> sl<33> vdd vss wl<67> / cell_PIM2
XI22739 bl<33> cbl<16> in1<66> in2<66> sl<33> vdd vss wl<66> / cell_PIM2
XI22737 bl<33> cbl<16> in1<69> in2<69> sl<33> vdd vss wl<69> / cell_PIM2
XI22736 bl<33> cbl<16> in1<68> in2<68> sl<33> vdd vss wl<68> / cell_PIM2
XI22088 bl<57> cbl<28> in1<93> in2<93> sl<57> vdd vss wl<93> / cell_PIM2
XI21434 bl<47> cbl<23> in1<108> in2<108> sl<47> vdd vss wl<108> / cell_PIM2
XI21433 bl<47> cbl<23> in1<109> in2<109> sl<47> vdd vss wl<109> / cell_PIM2
XI21432 bl<47> cbl<23> in1<110> in2<110> sl<47> vdd vss wl<110> / cell_PIM2
XI21431 bl<47> cbl<23> in1<111> in2<111> sl<47> vdd vss wl<111> / cell_PIM2
XI21430 bl<47> cbl<23> in1<112> in2<112> sl<47> vdd vss wl<112> / cell_PIM2
XI22082 bl<55> cbl<27> in1<89> in2<89> sl<55> vdd vss wl<89> / cell_PIM2
XI22081 bl<55> cbl<27> in1<90> in2<90> sl<55> vdd vss wl<90> / cell_PIM2
XI22080 bl<55> cbl<27> in1<91> in2<91> sl<55> vdd vss wl<91> / cell_PIM2
XI22079 bl<55> cbl<27> in1<92> in2<92> sl<55> vdd vss wl<92> / cell_PIM2
XI22730 bl<63> cbl<31> in1<70> in2<70> sl<63> vdd vss wl<70> / cell_PIM2
XI22729 bl<63> cbl<31> in1<71> in2<71> sl<63> vdd vss wl<71> / cell_PIM2
XI21424 bl<45> cbl<22> in1<110> in2<110> sl<45> vdd vss wl<110> / cell_PIM2
XI22078 bl<55> cbl<27> in1<93> in2<93> sl<55> vdd vss wl<93> / cell_PIM2
XI22727 bl<63> cbl<31> in1<73> in2<73> sl<63> vdd vss wl<73> / cell_PIM2
XI22726 bl<63> cbl<31> in1<74> in2<74> sl<63> vdd vss wl<74> / cell_PIM2
XI21423 bl<45> cbl<22> in1<109> in2<109> sl<45> vdd vss wl<109> / cell_PIM2
XI21422 bl<45> cbl<22> in1<108> in2<108> sl<45> vdd vss wl<108> / cell_PIM2
XI21421 bl<45> cbl<22> in1<112> in2<112> sl<45> vdd vss wl<112> / cell_PIM2
XI21420 bl<45> cbl<22> in1<111> in2<111> sl<45> vdd vss wl<111> / cell_PIM2
XI22072 bl<53> cbl<26> in1<91> in2<91> sl<53> vdd vss wl<91> / cell_PIM2
XI22071 bl<53> cbl<26> in1<90> in2<90> sl<53> vdd vss wl<90> / cell_PIM2
XI22070 bl<53> cbl<26> in1<89> in2<89> sl<53> vdd vss wl<89> / cell_PIM2
XI22069 bl<53> cbl<26> in1<93> in2<93> sl<53> vdd vss wl<93> / cell_PIM2
XI22720 bl<61> cbl<30> in1<71> in2<71> sl<61> vdd vss wl<71> / cell_PIM2
XI22719 bl<61> cbl<30> in1<70> in2<70> sl<61> vdd vss wl<70> / cell_PIM2
XI22717 bl<61> cbl<30> in1<73> in2<73> sl<61> vdd vss wl<73> / cell_PIM2
XI22716 bl<61> cbl<30> in1<72> in2<72> sl<61> vdd vss wl<72> / cell_PIM2
XI22068 bl<53> cbl<26> in1<92> in2<92> sl<53> vdd vss wl<92> / cell_PIM2
XI21414 bl<43> cbl<21> in1<108> in2<108> sl<43> vdd vss wl<108> / cell_PIM2
XI21413 bl<43> cbl<21> in1<109> in2<109> sl<43> vdd vss wl<109> / cell_PIM2
XI21412 bl<43> cbl<21> in1<110> in2<110> sl<43> vdd vss wl<110> / cell_PIM2
XI21411 bl<43> cbl<21> in1<111> in2<111> sl<43> vdd vss wl<111> / cell_PIM2
XI21410 bl<43> cbl<21> in1<112> in2<112> sl<43> vdd vss wl<112> / cell_PIM2
XI22062 bl<51> cbl<25> in1<89> in2<89> sl<51> vdd vss wl<89> / cell_PIM2
XI22061 bl<51> cbl<25> in1<90> in2<90> sl<51> vdd vss wl<90> / cell_PIM2
XI22060 bl<51> cbl<25> in1<91> in2<91> sl<51> vdd vss wl<91> / cell_PIM2
XI22059 bl<51> cbl<25> in1<92> in2<92> sl<51> vdd vss wl<92> / cell_PIM2
XI22710 bl<59> cbl<29> in1<70> in2<70> sl<59> vdd vss wl<70> / cell_PIM2
XI22709 bl<59> cbl<29> in1<71> in2<71> sl<59> vdd vss wl<71> / cell_PIM2
XI21404 bl<41> cbl<20> in1<108> in2<108> sl<41> vdd vss wl<108> / cell_PIM2
XI22058 bl<51> cbl<25> in1<93> in2<93> sl<51> vdd vss wl<93> / cell_PIM2
XI22707 bl<59> cbl<29> in1<73> in2<73> sl<59> vdd vss wl<73> / cell_PIM2
XI22706 bl<59> cbl<29> in1<74> in2<74> sl<59> vdd vss wl<74> / cell_PIM2
XI21403 bl<41> cbl<20> in1<109> in2<109> sl<41> vdd vss wl<109> / cell_PIM2
XI21402 bl<41> cbl<20> in1<110> in2<110> sl<41> vdd vss wl<110> / cell_PIM2
XI21401 bl<41> cbl<20> in1<111> in2<111> sl<41> vdd vss wl<111> / cell_PIM2
XI21400 bl<41> cbl<20> in1<112> in2<112> sl<41> vdd vss wl<112> / cell_PIM2
XI22052 bl<49> cbl<24> in1<91> in2<91> sl<49> vdd vss wl<91> / cell_PIM2
XI22051 bl<49> cbl<24> in1<90> in2<90> sl<49> vdd vss wl<90> / cell_PIM2
XI22050 bl<49> cbl<24> in1<89> in2<89> sl<49> vdd vss wl<89> / cell_PIM2
XI22049 bl<49> cbl<24> in1<93> in2<93> sl<49> vdd vss wl<93> / cell_PIM2
XI22700 bl<57> cbl<28> in1<70> in2<70> sl<57> vdd vss wl<70> / cell_PIM2
XI22699 bl<57> cbl<28> in1<71> in2<71> sl<57> vdd vss wl<71> / cell_PIM2
XI22697 bl<57> cbl<28> in1<73> in2<73> sl<57> vdd vss wl<73> / cell_PIM2
XI22696 bl<57> cbl<28> in1<74> in2<74> sl<57> vdd vss wl<74> / cell_PIM2
XI22048 bl<49> cbl<24> in1<92> in2<92> sl<49> vdd vss wl<92> / cell_PIM2
XI21394 bl<39> cbl<19> in1<108> in2<108> sl<39> vdd vss wl<108> / cell_PIM2
XI21393 bl<39> cbl<19> in1<109> in2<109> sl<39> vdd vss wl<109> / cell_PIM2
XI21392 bl<39> cbl<19> in1<110> in2<110> sl<39> vdd vss wl<110> / cell_PIM2
XI21391 bl<39> cbl<19> in1<111> in2<111> sl<39> vdd vss wl<111> / cell_PIM2
XI21390 bl<39> cbl<19> in1<112> in2<112> sl<39> vdd vss wl<112> / cell_PIM2
XI22042 bl<47> cbl<23> in1<89> in2<89> sl<47> vdd vss wl<89> / cell_PIM2
XI22041 bl<47> cbl<23> in1<90> in2<90> sl<47> vdd vss wl<90> / cell_PIM2
XI22040 bl<47> cbl<23> in1<91> in2<91> sl<47> vdd vss wl<91> / cell_PIM2
XI22039 bl<47> cbl<23> in1<92> in2<92> sl<47> vdd vss wl<92> / cell_PIM2
XI22690 bl<55> cbl<27> in1<70> in2<70> sl<55> vdd vss wl<70> / cell_PIM2
XI22689 bl<55> cbl<27> in1<71> in2<71> sl<55> vdd vss wl<71> / cell_PIM2
XI21384 bl<37> cbl<18> in1<110> in2<110> sl<37> vdd vss wl<110> / cell_PIM2
XI22038 bl<47> cbl<23> in1<93> in2<93> sl<47> vdd vss wl<93> / cell_PIM2
XI22687 bl<55> cbl<27> in1<73> in2<73> sl<55> vdd vss wl<73> / cell_PIM2
XI22686 bl<55> cbl<27> in1<74> in2<74> sl<55> vdd vss wl<74> / cell_PIM2
XI21383 bl<37> cbl<18> in1<109> in2<109> sl<37> vdd vss wl<109> / cell_PIM2
XI21382 bl<37> cbl<18> in1<108> in2<108> sl<37> vdd vss wl<108> / cell_PIM2
XI21381 bl<37> cbl<18> in1<112> in2<112> sl<37> vdd vss wl<112> / cell_PIM2
XI21380 bl<37> cbl<18> in1<111> in2<111> sl<37> vdd vss wl<111> / cell_PIM2
XI22032 bl<45> cbl<22> in1<91> in2<91> sl<45> vdd vss wl<91> / cell_PIM2
XI22031 bl<45> cbl<22> in1<90> in2<90> sl<45> vdd vss wl<90> / cell_PIM2
XI22030 bl<45> cbl<22> in1<89> in2<89> sl<45> vdd vss wl<89> / cell_PIM2
XI22029 bl<45> cbl<22> in1<93> in2<93> sl<45> vdd vss wl<93> / cell_PIM2
XI22680 bl<53> cbl<26> in1<71> in2<71> sl<53> vdd vss wl<71> / cell_PIM2
XI22679 bl<53> cbl<26> in1<70> in2<70> sl<53> vdd vss wl<70> / cell_PIM2
XI22677 bl<53> cbl<26> in1<73> in2<73> sl<53> vdd vss wl<73> / cell_PIM2
XI22676 bl<53> cbl<26> in1<72> in2<72> sl<53> vdd vss wl<72> / cell_PIM2
XI22028 bl<45> cbl<22> in1<92> in2<92> sl<45> vdd vss wl<92> / cell_PIM2
XI21374 bl<35> cbl<17> in1<108> in2<108> sl<35> vdd vss wl<108> / cell_PIM2
XI21373 bl<35> cbl<17> in1<109> in2<109> sl<35> vdd vss wl<109> / cell_PIM2
XI21372 bl<35> cbl<17> in1<110> in2<110> sl<35> vdd vss wl<110> / cell_PIM2
XI21371 bl<35> cbl<17> in1<111> in2<111> sl<35> vdd vss wl<111> / cell_PIM2
XI21370 bl<35> cbl<17> in1<112> in2<112> sl<35> vdd vss wl<112> / cell_PIM2
XI22022 bl<43> cbl<21> in1<89> in2<89> sl<43> vdd vss wl<89> / cell_PIM2
XI22021 bl<43> cbl<21> in1<90> in2<90> sl<43> vdd vss wl<90> / cell_PIM2
XI22020 bl<43> cbl<21> in1<91> in2<91> sl<43> vdd vss wl<91> / cell_PIM2
XI22019 bl<43> cbl<21> in1<92> in2<92> sl<43> vdd vss wl<92> / cell_PIM2
XI22670 bl<51> cbl<25> in1<70> in2<70> sl<51> vdd vss wl<70> / cell_PIM2
XI22669 bl<51> cbl<25> in1<71> in2<71> sl<51> vdd vss wl<71> / cell_PIM2
XI21364 bl<33> cbl<16> in1<110> in2<110> sl<33> vdd vss wl<110> / cell_PIM2
XI22018 bl<43> cbl<21> in1<93> in2<93> sl<43> vdd vss wl<93> / cell_PIM2
XI22667 bl<51> cbl<25> in1<73> in2<73> sl<51> vdd vss wl<73> / cell_PIM2
XI22666 bl<51> cbl<25> in1<74> in2<74> sl<51> vdd vss wl<74> / cell_PIM2
XI21363 bl<33> cbl<16> in1<109> in2<109> sl<33> vdd vss wl<109> / cell_PIM2
XI21362 bl<33> cbl<16> in1<108> in2<108> sl<33> vdd vss wl<108> / cell_PIM2
XI21361 bl<33> cbl<16> in1<112> in2<112> sl<33> vdd vss wl<112> / cell_PIM2
XI21360 bl<33> cbl<16> in1<111> in2<111> sl<33> vdd vss wl<111> / cell_PIM2
XI22012 bl<41> cbl<20> in1<89> in2<89> sl<41> vdd vss wl<89> / cell_PIM2
XI22011 bl<41> cbl<20> in1<90> in2<90> sl<41> vdd vss wl<90> / cell_PIM2
XI22010 bl<41> cbl<20> in1<91> in2<91> sl<41> vdd vss wl<91> / cell_PIM2
XI22009 bl<41> cbl<20> in1<92> in2<92> sl<41> vdd vss wl<92> / cell_PIM2
XI22660 bl<49> cbl<24> in1<71> in2<71> sl<49> vdd vss wl<71> / cell_PIM2
XI22659 bl<49> cbl<24> in1<70> in2<70> sl<49> vdd vss wl<70> / cell_PIM2
XI22657 bl<49> cbl<24> in1<73> in2<73> sl<49> vdd vss wl<73> / cell_PIM2
XI22656 bl<49> cbl<24> in1<72> in2<72> sl<49> vdd vss wl<72> / cell_PIM2
XI22008 bl<41> cbl<20> in1<93> in2<93> sl<41> vdd vss wl<93> / cell_PIM2
XI21354 bl<63> cbl<31> in1<113> in2<113> sl<63> vdd vss wl<113> / cell_PIM2
XI21353 bl<63> cbl<31> in1<114> in2<114> sl<63> vdd vss wl<114> / cell_PIM2
XI21352 bl<63> cbl<31> in1<115> in2<115> sl<63> vdd vss wl<115> / cell_PIM2
XI21351 bl<63> cbl<31> in1<116> in2<116> sl<63> vdd vss wl<116> / cell_PIM2
XI21350 bl<63> cbl<31> in1<117> in2<117> sl<63> vdd vss wl<117> / cell_PIM2
XI22002 bl<39> cbl<19> in1<89> in2<89> sl<39> vdd vss wl<89> / cell_PIM2
XI22001 bl<39> cbl<19> in1<90> in2<90> sl<39> vdd vss wl<90> / cell_PIM2
XI22000 bl<39> cbl<19> in1<91> in2<91> sl<39> vdd vss wl<91> / cell_PIM2
XI21999 bl<39> cbl<19> in1<92> in2<92> sl<39> vdd vss wl<92> / cell_PIM2
XI22650 bl<47> cbl<23> in1<70> in2<70> sl<47> vdd vss wl<70> / cell_PIM2
XI22649 bl<47> cbl<23> in1<71> in2<71> sl<47> vdd vss wl<71> / cell_PIM2
XI21344 bl<61> cbl<30> in1<115> in2<115> sl<61> vdd vss wl<115> / cell_PIM2
XI21998 bl<39> cbl<19> in1<93> in2<93> sl<39> vdd vss wl<93> / cell_PIM2
XI22647 bl<47> cbl<23> in1<73> in2<73> sl<47> vdd vss wl<73> / cell_PIM2
XI22646 bl<47> cbl<23> in1<74> in2<74> sl<47> vdd vss wl<74> / cell_PIM2
XI21343 bl<61> cbl<30> in1<114> in2<114> sl<61> vdd vss wl<114> / cell_PIM2
XI21342 bl<61> cbl<30> in1<113> in2<113> sl<61> vdd vss wl<113> / cell_PIM2
XI21341 bl<61> cbl<30> in1<117> in2<117> sl<61> vdd vss wl<117> / cell_PIM2
XI21340 bl<61> cbl<30> in1<116> in2<116> sl<61> vdd vss wl<116> / cell_PIM2
XI21992 bl<37> cbl<18> in1<91> in2<91> sl<37> vdd vss wl<91> / cell_PIM2
XI21991 bl<37> cbl<18> in1<90> in2<90> sl<37> vdd vss wl<90> / cell_PIM2
XI21990 bl<37> cbl<18> in1<89> in2<89> sl<37> vdd vss wl<89> / cell_PIM2
XI21989 bl<37> cbl<18> in1<93> in2<93> sl<37> vdd vss wl<93> / cell_PIM2
XI22640 bl<45> cbl<22> in1<71> in2<71> sl<45> vdd vss wl<71> / cell_PIM2
XI22639 bl<45> cbl<22> in1<70> in2<70> sl<45> vdd vss wl<70> / cell_PIM2
XI22637 bl<45> cbl<22> in1<73> in2<73> sl<45> vdd vss wl<73> / cell_PIM2
XI22636 bl<45> cbl<22> in1<72> in2<72> sl<45> vdd vss wl<72> / cell_PIM2
XI21988 bl<37> cbl<18> in1<92> in2<92> sl<37> vdd vss wl<92> / cell_PIM2
XI21334 bl<59> cbl<29> in1<113> in2<113> sl<59> vdd vss wl<113> / cell_PIM2
XI21333 bl<59> cbl<29> in1<114> in2<114> sl<59> vdd vss wl<114> / cell_PIM2
XI21332 bl<59> cbl<29> in1<115> in2<115> sl<59> vdd vss wl<115> / cell_PIM2
XI21331 bl<59> cbl<29> in1<116> in2<116> sl<59> vdd vss wl<116> / cell_PIM2
XI21330 bl<59> cbl<29> in1<117> in2<117> sl<59> vdd vss wl<117> / cell_PIM2
XI21982 bl<35> cbl<17> in1<89> in2<89> sl<35> vdd vss wl<89> / cell_PIM2
XI21981 bl<35> cbl<17> in1<90> in2<90> sl<35> vdd vss wl<90> / cell_PIM2
XI21980 bl<35> cbl<17> in1<91> in2<91> sl<35> vdd vss wl<91> / cell_PIM2
XI21979 bl<35> cbl<17> in1<92> in2<92> sl<35> vdd vss wl<92> / cell_PIM2
XI22630 bl<43> cbl<21> in1<70> in2<70> sl<43> vdd vss wl<70> / cell_PIM2
XI22629 bl<43> cbl<21> in1<71> in2<71> sl<43> vdd vss wl<71> / cell_PIM2
XI21324 bl<57> cbl<28> in1<113> in2<113> sl<57> vdd vss wl<113> / cell_PIM2
XI21978 bl<35> cbl<17> in1<93> in2<93> sl<35> vdd vss wl<93> / cell_PIM2
XI22627 bl<43> cbl<21> in1<73> in2<73> sl<43> vdd vss wl<73> / cell_PIM2
XI22626 bl<43> cbl<21> in1<74> in2<74> sl<43> vdd vss wl<74> / cell_PIM2
XI21323 bl<57> cbl<28> in1<114> in2<114> sl<57> vdd vss wl<114> / cell_PIM2
XI21322 bl<57> cbl<28> in1<115> in2<115> sl<57> vdd vss wl<115> / cell_PIM2
XI21321 bl<57> cbl<28> in1<116> in2<116> sl<57> vdd vss wl<116> / cell_PIM2
XI21320 bl<57> cbl<28> in1<117> in2<117> sl<57> vdd vss wl<117> / cell_PIM2
XI21972 bl<33> cbl<16> in1<91> in2<91> sl<33> vdd vss wl<91> / cell_PIM2
XI21971 bl<33> cbl<16> in1<90> in2<90> sl<33> vdd vss wl<90> / cell_PIM2
XI21970 bl<33> cbl<16> in1<89> in2<89> sl<33> vdd vss wl<89> / cell_PIM2
XI21969 bl<33> cbl<16> in1<93> in2<93> sl<33> vdd vss wl<93> / cell_PIM2
XI22620 bl<41> cbl<20> in1<70> in2<70> sl<41> vdd vss wl<70> / cell_PIM2
XI22619 bl<41> cbl<20> in1<71> in2<71> sl<41> vdd vss wl<71> / cell_PIM2
XI22617 bl<41> cbl<20> in1<73> in2<73> sl<41> vdd vss wl<73> / cell_PIM2
XI22616 bl<41> cbl<20> in1<74> in2<74> sl<41> vdd vss wl<74> / cell_PIM2
XI21968 bl<33> cbl<16> in1<92> in2<92> sl<33> vdd vss wl<92> / cell_PIM2
XI21314 bl<55> cbl<27> in1<113> in2<113> sl<55> vdd vss wl<113> / cell_PIM2
XI21313 bl<55> cbl<27> in1<114> in2<114> sl<55> vdd vss wl<114> / cell_PIM2
XI21312 bl<55> cbl<27> in1<115> in2<115> sl<55> vdd vss wl<115> / cell_PIM2
XI21311 bl<55> cbl<27> in1<116> in2<116> sl<55> vdd vss wl<116> / cell_PIM2
XI21310 bl<55> cbl<27> in1<117> in2<117> sl<55> vdd vss wl<117> / cell_PIM2
XI21962 bl<63> cbl<31> in1<94> in2<94> sl<63> vdd vss wl<94> / cell_PIM2
XI21961 bl<63> cbl<31> in1<95> in2<95> sl<63> vdd vss wl<95> / cell_PIM2
XI21960 bl<63> cbl<31> in1<96> in2<96> sl<63> vdd vss wl<96> / cell_PIM2
XI21959 bl<63> cbl<31> in1<97> in2<97> sl<63> vdd vss wl<97> / cell_PIM2
XI22610 bl<39> cbl<19> in1<70> in2<70> sl<39> vdd vss wl<70> / cell_PIM2
XI22609 bl<39> cbl<19> in1<71> in2<71> sl<39> vdd vss wl<71> / cell_PIM2
XI21304 bl<53> cbl<26> in1<115> in2<115> sl<53> vdd vss wl<115> / cell_PIM2
XI21958 bl<63> cbl<31> in1<98> in2<98> sl<63> vdd vss wl<98> / cell_PIM2
XI22607 bl<39> cbl<19> in1<73> in2<73> sl<39> vdd vss wl<73> / cell_PIM2
XI22606 bl<39> cbl<19> in1<74> in2<74> sl<39> vdd vss wl<74> / cell_PIM2
XI21303 bl<53> cbl<26> in1<114> in2<114> sl<53> vdd vss wl<114> / cell_PIM2
XI21302 bl<53> cbl<26> in1<113> in2<113> sl<53> vdd vss wl<113> / cell_PIM2
XI21301 bl<53> cbl<26> in1<117> in2<117> sl<53> vdd vss wl<117> / cell_PIM2
XI21300 bl<53> cbl<26> in1<116> in2<116> sl<53> vdd vss wl<116> / cell_PIM2
XI21952 bl<61> cbl<30> in1<95> in2<95> sl<61> vdd vss wl<95> / cell_PIM2
XI21951 bl<61> cbl<30> in1<94> in2<94> sl<61> vdd vss wl<94> / cell_PIM2
XI21950 bl<61> cbl<30> in1<98> in2<98> sl<61> vdd vss wl<98> / cell_PIM2
XI21949 bl<61> cbl<30> in1<97> in2<97> sl<61> vdd vss wl<97> / cell_PIM2
XI22600 bl<37> cbl<18> in1<71> in2<71> sl<37> vdd vss wl<71> / cell_PIM2
XI22599 bl<37> cbl<18> in1<70> in2<70> sl<37> vdd vss wl<70> / cell_PIM2
XI22597 bl<37> cbl<18> in1<73> in2<73> sl<37> vdd vss wl<73> / cell_PIM2
XI22596 bl<37> cbl<18> in1<72> in2<72> sl<37> vdd vss wl<72> / cell_PIM2
XI21948 bl<61> cbl<30> in1<96> in2<96> sl<61> vdd vss wl<96> / cell_PIM2
XI21294 bl<51> cbl<25> in1<113> in2<113> sl<51> vdd vss wl<113> / cell_PIM2
XI21293 bl<51> cbl<25> in1<114> in2<114> sl<51> vdd vss wl<114> / cell_PIM2
XI21292 bl<51> cbl<25> in1<115> in2<115> sl<51> vdd vss wl<115> / cell_PIM2
XI21291 bl<51> cbl<25> in1<116> in2<116> sl<51> vdd vss wl<116> / cell_PIM2
XI21290 bl<51> cbl<25> in1<117> in2<117> sl<51> vdd vss wl<117> / cell_PIM2
XI21942 bl<59> cbl<29> in1<94> in2<94> sl<59> vdd vss wl<94> / cell_PIM2
XI21941 bl<59> cbl<29> in1<95> in2<95> sl<59> vdd vss wl<95> / cell_PIM2
XI21940 bl<59> cbl<29> in1<96> in2<96> sl<59> vdd vss wl<96> / cell_PIM2
XI21939 bl<59> cbl<29> in1<97> in2<97> sl<59> vdd vss wl<97> / cell_PIM2
XI22590 bl<35> cbl<17> in1<70> in2<70> sl<35> vdd vss wl<70> / cell_PIM2
XI22589 bl<35> cbl<17> in1<71> in2<71> sl<35> vdd vss wl<71> / cell_PIM2
XI21284 bl<49> cbl<24> in1<115> in2<115> sl<49> vdd vss wl<115> / cell_PIM2
XI21938 bl<59> cbl<29> in1<98> in2<98> sl<59> vdd vss wl<98> / cell_PIM2
XI22587 bl<35> cbl<17> in1<73> in2<73> sl<35> vdd vss wl<73> / cell_PIM2
XI22586 bl<35> cbl<17> in1<74> in2<74> sl<35> vdd vss wl<74> / cell_PIM2
XI21283 bl<49> cbl<24> in1<114> in2<114> sl<49> vdd vss wl<114> / cell_PIM2
XI21282 bl<49> cbl<24> in1<113> in2<113> sl<49> vdd vss wl<113> / cell_PIM2
XI21281 bl<49> cbl<24> in1<117> in2<117> sl<49> vdd vss wl<117> / cell_PIM2
XI21280 bl<49> cbl<24> in1<116> in2<116> sl<49> vdd vss wl<116> / cell_PIM2
XI21932 bl<57> cbl<28> in1<94> in2<94> sl<57> vdd vss wl<94> / cell_PIM2
XI21931 bl<57> cbl<28> in1<95> in2<95> sl<57> vdd vss wl<95> / cell_PIM2
XI21930 bl<57> cbl<28> in1<96> in2<96> sl<57> vdd vss wl<96> / cell_PIM2
XI21929 bl<57> cbl<28> in1<97> in2<97> sl<57> vdd vss wl<97> / cell_PIM2
XI22580 bl<33> cbl<16> in1<71> in2<71> sl<33> vdd vss wl<71> / cell_PIM2
XI22579 bl<33> cbl<16> in1<70> in2<70> sl<33> vdd vss wl<70> / cell_PIM2
XI22577 bl<33> cbl<16> in1<73> in2<73> sl<33> vdd vss wl<73> / cell_PIM2
XI22576 bl<33> cbl<16> in1<72> in2<72> sl<33> vdd vss wl<72> / cell_PIM2
XI21928 bl<57> cbl<28> in1<98> in2<98> sl<57> vdd vss wl<98> / cell_PIM2
XI21274 bl<47> cbl<23> in1<113> in2<113> sl<47> vdd vss wl<113> / cell_PIM2
XI21273 bl<47> cbl<23> in1<114> in2<114> sl<47> vdd vss wl<114> / cell_PIM2
XI21272 bl<47> cbl<23> in1<115> in2<115> sl<47> vdd vss wl<115> / cell_PIM2
XI21271 bl<47> cbl<23> in1<116> in2<116> sl<47> vdd vss wl<116> / cell_PIM2
XI21270 bl<47> cbl<23> in1<117> in2<117> sl<47> vdd vss wl<117> / cell_PIM2
XI21922 bl<55> cbl<27> in1<94> in2<94> sl<55> vdd vss wl<94> / cell_PIM2
XI21921 bl<55> cbl<27> in1<95> in2<95> sl<55> vdd vss wl<95> / cell_PIM2
XI21920 bl<55> cbl<27> in1<96> in2<96> sl<55> vdd vss wl<96> / cell_PIM2
XI21919 bl<55> cbl<27> in1<97> in2<97> sl<55> vdd vss wl<97> / cell_PIM2
XI22570 bl<63> cbl<31> in1<75> in2<75> sl<63> vdd vss wl<75> / cell_PIM2
XI22569 bl<63> cbl<31> in1<76> in2<76> sl<63> vdd vss wl<76> / cell_PIM2
XI21264 bl<45> cbl<22> in1<115> in2<115> sl<45> vdd vss wl<115> / cell_PIM2
XI21918 bl<55> cbl<27> in1<98> in2<98> sl<55> vdd vss wl<98> / cell_PIM2
XI22567 bl<63> cbl<31> in1<78> in2<78> sl<63> vdd vss wl<78> / cell_PIM2
XI22566 bl<63> cbl<31> in1<79> in2<79> sl<63> vdd vss wl<79> / cell_PIM2
XI19762 bl<17> cbl<8> in1<65> in2<65> sl<17> vdd vss wl<65> / cell_PIM2
XI19761 bl<17> cbl<8> in1<69> in2<69> sl<17> vdd vss wl<69> / cell_PIM2
XI19760 bl<17> cbl<8> in1<68> in2<68> sl<17> vdd vss wl<68> / cell_PIM2
XI19763 bl<17> cbl<8> in1<66> in2<66> sl<17> vdd vss wl<66> / cell_PIM2
XI20282 bl<31> cbl<15> in1<37> in2<37> sl<31> vdd vss wl<37> / cell_PIM2
XI20281 bl<31> cbl<15> in1<38> in2<38> sl<31> vdd vss wl<38> / cell_PIM2
XI20933 bl<43> cbl<21> in1<126> in2<126> sl<43> vdd vss wl<126> / cell_PIM2
XI20932 bl<43> cbl<21> in1<125> in2<125> sl<43> vdd vss wl<125> / cell_PIM2
XI20931 bl<43> cbl<21> in1<123> in2<123> sl<43> vdd vss wl<123> / cell_PIM2
XI20930 bl<43> cbl<21> in1<124> in2<124> sl<43> vdd vss wl<124> / cell_PIM2
XI20924 bl<41> cbl<20> in1<127> in2<127> sl<41> vdd vss wl<127> / cell_PIM2
XI20280 bl<31> cbl<15> in1<39> in2<39> sl<31> vdd vss wl<39> / cell_PIM2
XI20279 bl<31> cbl<15> in1<40> in2<40> sl<31> vdd vss wl<40> / cell_PIM2
XI19754 bl<31> cbl<15> in1<70> in2<70> sl<31> vdd vss wl<70> / cell_PIM2
XI19752 bl<31> cbl<15> in1<72> in2<72> sl<31> vdd vss wl<72> / cell_PIM2
XI19751 bl<31> cbl<15> in1<73> in2<73> sl<31> vdd vss wl<73> / cell_PIM2
XI19750 bl<31> cbl<15> in1<74> in2<74> sl<31> vdd vss wl<74> / cell_PIM2
XI19753 bl<31> cbl<15> in1<71> in2<71> sl<31> vdd vss wl<71> / cell_PIM2
XI20274 bl<29> cbl<14> in1<38> in2<38> sl<29> vdd vss wl<38> / cell_PIM2
XI20273 bl<29> cbl<14> in1<37> in2<37> sl<29> vdd vss wl<37> / cell_PIM2
XI20923 bl<41> cbl<20> in1<126> in2<126> sl<41> vdd vss wl<126> / cell_PIM2
XI20922 bl<41> cbl<20> in1<125> in2<125> sl<41> vdd vss wl<125> / cell_PIM2
XI20921 bl<41> cbl<20> in1<123> in2<123> sl<41> vdd vss wl<123> / cell_PIM2
XI20920 bl<41> cbl<20> in1<124> in2<124> sl<41> vdd vss wl<124> / cell_PIM2
XI19744 bl<29> cbl<14> in1<71> in2<71> sl<29> vdd vss wl<71> / cell_PIM2
XI20272 bl<29> cbl<14> in1<40> in2<40> sl<29> vdd vss wl<40> / cell_PIM2
XI20271 bl<29> cbl<14> in1<39> in2<39> sl<29> vdd vss wl<39> / cell_PIM2
XI20914 bl<39> cbl<19> in1<127> in2<127> sl<39> vdd vss wl<127> / cell_PIM2
XI19742 bl<29> cbl<14> in1<74> in2<74> sl<29> vdd vss wl<74> / cell_PIM2
XI19741 bl<29> cbl<14> in1<73> in2<73> sl<29> vdd vss wl<73> / cell_PIM2
XI19740 bl<29> cbl<14> in1<72> in2<72> sl<29> vdd vss wl<72> / cell_PIM2
XI19743 bl<29> cbl<14> in1<70> in2<70> sl<29> vdd vss wl<70> / cell_PIM2
XI20266 bl<27> cbl<13> in1<37> in2<37> sl<27> vdd vss wl<37> / cell_PIM2
XI20265 bl<27> cbl<13> in1<38> in2<38> sl<27> vdd vss wl<38> / cell_PIM2
XI20913 bl<39> cbl<19> in1<126> in2<126> sl<39> vdd vss wl<126> / cell_PIM2
XI20912 bl<39> cbl<19> in1<125> in2<125> sl<39> vdd vss wl<125> / cell_PIM2
XI20911 bl<39> cbl<19> in1<123> in2<123> sl<39> vdd vss wl<123> / cell_PIM2
XI20910 bl<39> cbl<19> in1<124> in2<124> sl<39> vdd vss wl<124> / cell_PIM2
XI20904 bl<37> cbl<18> in1<127> in2<127> sl<37> vdd vss wl<127> / cell_PIM2
XI20264 bl<27> cbl<13> in1<39> in2<39> sl<27> vdd vss wl<39> / cell_PIM2
XI20263 bl<27> cbl<13> in1<40> in2<40> sl<27> vdd vss wl<40> / cell_PIM2
XI19734 bl<27> cbl<13> in1<70> in2<70> sl<27> vdd vss wl<70> / cell_PIM2
XI19732 bl<27> cbl<13> in1<72> in2<72> sl<27> vdd vss wl<72> / cell_PIM2
XI19731 bl<27> cbl<13> in1<73> in2<73> sl<27> vdd vss wl<73> / cell_PIM2
XI19730 bl<27> cbl<13> in1<74> in2<74> sl<27> vdd vss wl<74> / cell_PIM2
XI19733 bl<27> cbl<13> in1<71> in2<71> sl<27> vdd vss wl<71> / cell_PIM2
XI20258 bl<25> cbl<12> in1<37> in2<37> sl<25> vdd vss wl<37> / cell_PIM2
XI20257 bl<25> cbl<12> in1<38> in2<38> sl<25> vdd vss wl<38> / cell_PIM2
XI20903 bl<37> cbl<18> in1<126> in2<126> sl<37> vdd vss wl<126> / cell_PIM2
XI20902 bl<37> cbl<18> in1<125> in2<125> sl<37> vdd vss wl<125> / cell_PIM2
XI20901 bl<37> cbl<18> in1<124> in2<124> sl<37> vdd vss wl<124> / cell_PIM2
XI20900 bl<37> cbl<18> in1<123> in2<123> sl<37> vdd vss wl<123> / cell_PIM2
XI19724 bl<25> cbl<12> in1<70> in2<70> sl<25> vdd vss wl<70> / cell_PIM2
XI20256 bl<25> cbl<12> in1<39> in2<39> sl<25> vdd vss wl<39> / cell_PIM2
XI20255 bl<25> cbl<12> in1<40> in2<40> sl<25> vdd vss wl<40> / cell_PIM2
XI20894 bl<35> cbl<17> in1<127> in2<127> sl<35> vdd vss wl<127> / cell_PIM2
XI19722 bl<25> cbl<12> in1<72> in2<72> sl<25> vdd vss wl<72> / cell_PIM2
XI19721 bl<25> cbl<12> in1<73> in2<73> sl<25> vdd vss wl<73> / cell_PIM2
XI19720 bl<25> cbl<12> in1<74> in2<74> sl<25> vdd vss wl<74> / cell_PIM2
XI19723 bl<25> cbl<12> in1<71> in2<71> sl<25> vdd vss wl<71> / cell_PIM2
XI20250 bl<23> cbl<11> in1<37> in2<37> sl<23> vdd vss wl<37> / cell_PIM2
XI20249 bl<23> cbl<11> in1<38> in2<38> sl<23> vdd vss wl<38> / cell_PIM2
XI20893 bl<35> cbl<17> in1<126> in2<126> sl<35> vdd vss wl<126> / cell_PIM2
XI20892 bl<35> cbl<17> in1<125> in2<125> sl<35> vdd vss wl<125> / cell_PIM2
XI20891 bl<35> cbl<17> in1<123> in2<123> sl<35> vdd vss wl<123> / cell_PIM2
XI20890 bl<35> cbl<17> in1<124> in2<124> sl<35> vdd vss wl<124> / cell_PIM2
XI20884 bl<33> cbl<16> in1<127> in2<127> sl<33> vdd vss wl<127> / cell_PIM2
XI20248 bl<23> cbl<11> in1<39> in2<39> sl<23> vdd vss wl<39> / cell_PIM2
XI20247 bl<23> cbl<11> in1<40> in2<40> sl<23> vdd vss wl<40> / cell_PIM2
XI19714 bl<23> cbl<11> in1<70> in2<70> sl<23> vdd vss wl<70> / cell_PIM2
XI19712 bl<23> cbl<11> in1<72> in2<72> sl<23> vdd vss wl<72> / cell_PIM2
XI19711 bl<23> cbl<11> in1<73> in2<73> sl<23> vdd vss wl<73> / cell_PIM2
XI19710 bl<23> cbl<11> in1<74> in2<74> sl<23> vdd vss wl<74> / cell_PIM2
XI19713 bl<23> cbl<11> in1<71> in2<71> sl<23> vdd vss wl<71> / cell_PIM2
XI20242 bl<21> cbl<10> in1<38> in2<38> sl<21> vdd vss wl<38> / cell_PIM2
XI20241 bl<21> cbl<10> in1<37> in2<37> sl<21> vdd vss wl<37> / cell_PIM2
XI20883 bl<33> cbl<16> in1<126> in2<126> sl<33> vdd vss wl<126> / cell_PIM2
XI20882 bl<33> cbl<16> in1<125> in2<125> sl<33> vdd vss wl<125> / cell_PIM2
XI20881 bl<33> cbl<16> in1<124> in2<124> sl<33> vdd vss wl<124> / cell_PIM2
XI20880 bl<33> cbl<16> in1<123> in2<123> sl<33> vdd vss wl<123> / cell_PIM2
XI19704 bl<21> cbl<10> in1<71> in2<71> sl<21> vdd vss wl<71> / cell_PIM2
XI20240 bl<21> cbl<10> in1<40> in2<40> sl<21> vdd vss wl<40> / cell_PIM2
XI20239 bl<21> cbl<10> in1<39> in2<39> sl<21> vdd vss wl<39> / cell_PIM2
XI20874 bl<31> cbl<15> in1<0> in2<0> sl<31> vdd vss wl<0> / cell_PIM2
XI19702 bl<21> cbl<10> in1<74> in2<74> sl<21> vdd vss wl<74> / cell_PIM2
XI19701 bl<21> cbl<10> in1<73> in2<73> sl<21> vdd vss wl<73> / cell_PIM2
XI19700 bl<21> cbl<10> in1<72> in2<72> sl<21> vdd vss wl<72> / cell_PIM2
XI19703 bl<21> cbl<10> in1<70> in2<70> sl<21> vdd vss wl<70> / cell_PIM2
XI20234 bl<19> cbl<9> in1<37> in2<37> sl<19> vdd vss wl<37> / cell_PIM2
XI20233 bl<19> cbl<9> in1<38> in2<38> sl<19> vdd vss wl<38> / cell_PIM2
XI20873 bl<31> cbl<15> in1<1> in2<1> sl<31> vdd vss wl<1> / cell_PIM2
XI20872 bl<31> cbl<15> in1<2> in2<2> sl<31> vdd vss wl<2> / cell_PIM2
XI20868 bl<29> cbl<14> in1<0> in2<0> sl<29> vdd vss wl<0> / cell_PIM2
XI20867 bl<29> cbl<14> in1<2> in2<2> sl<29> vdd vss wl<2> / cell_PIM2
XI20866 bl<29> cbl<14> in1<1> in2<1> sl<29> vdd vss wl<1> / cell_PIM2
XI20232 bl<19> cbl<9> in1<39> in2<39> sl<19> vdd vss wl<39> / cell_PIM2
XI20231 bl<19> cbl<9> in1<40> in2<40> sl<19> vdd vss wl<40> / cell_PIM2
XI19694 bl<19> cbl<9> in1<70> in2<70> sl<19> vdd vss wl<70> / cell_PIM2
XI19692 bl<19> cbl<9> in1<72> in2<72> sl<19> vdd vss wl<72> / cell_PIM2
XI19691 bl<19> cbl<9> in1<73> in2<73> sl<19> vdd vss wl<73> / cell_PIM2
XI19690 bl<19> cbl<9> in1<74> in2<74> sl<19> vdd vss wl<74> / cell_PIM2
XI19693 bl<19> cbl<9> in1<71> in2<71> sl<19> vdd vss wl<71> / cell_PIM2
XI20226 bl<17> cbl<8> in1<38> in2<38> sl<17> vdd vss wl<38> / cell_PIM2
XI20225 bl<17> cbl<8> in1<37> in2<37> sl<17> vdd vss wl<37> / cell_PIM2
XI20862 bl<27> cbl<13> in1<0> in2<0> sl<27> vdd vss wl<0> / cell_PIM2
XI20861 bl<27> cbl<13> in1<1> in2<1> sl<27> vdd vss wl<1> / cell_PIM2
XI20860 bl<27> cbl<13> in1<2> in2<2> sl<27> vdd vss wl<2> / cell_PIM2
XI19684 bl<17> cbl<8> in1<71> in2<71> sl<17> vdd vss wl<71> / cell_PIM2
XI20224 bl<17> cbl<8> in1<40> in2<40> sl<17> vdd vss wl<40> / cell_PIM2
XI20223 bl<17> cbl<8> in1<39> in2<39> sl<17> vdd vss wl<39> / cell_PIM2
XI20856 bl<25> cbl<12> in1<0> in2<0> sl<25> vdd vss wl<0> / cell_PIM2
XI20855 bl<25> cbl<12> in1<1> in2<1> sl<25> vdd vss wl<1> / cell_PIM2
XI20854 bl<25> cbl<12> in1<2> in2<2> sl<25> vdd vss wl<2> / cell_PIM2
XI19682 bl<17> cbl<8> in1<74> in2<74> sl<17> vdd vss wl<74> / cell_PIM2
XI19681 bl<17> cbl<8> in1<73> in2<73> sl<17> vdd vss wl<73> / cell_PIM2
XI19680 bl<17> cbl<8> in1<72> in2<72> sl<17> vdd vss wl<72> / cell_PIM2
XI19683 bl<17> cbl<8> in1<70> in2<70> sl<17> vdd vss wl<70> / cell_PIM2
XI20218 bl<31> cbl<15> in1<41> in2<41> sl<31> vdd vss wl<41> / cell_PIM2
XI20217 bl<31> cbl<15> in1<42> in2<42> sl<31> vdd vss wl<42> / cell_PIM2
XI20850 bl<23> cbl<11> in1<0> in2<0> sl<23> vdd vss wl<0> / cell_PIM2
XI20849 bl<23> cbl<11> in1<1> in2<1> sl<23> vdd vss wl<1> / cell_PIM2
XI20848 bl<23> cbl<11> in1<2> in2<2> sl<23> vdd vss wl<2> / cell_PIM2
XI20844 bl<21> cbl<10> in1<0> in2<0> sl<21> vdd vss wl<0> / cell_PIM2
XI20216 bl<31> cbl<15> in1<43> in2<43> sl<31> vdd vss wl<43> / cell_PIM2
XI20215 bl<31> cbl<15> in1<44> in2<44> sl<31> vdd vss wl<44> / cell_PIM2
XI20214 bl<31> cbl<15> in1<45> in2<45> sl<31> vdd vss wl<45> / cell_PIM2
XI19674 bl<31> cbl<15> in1<75> in2<75> sl<31> vdd vss wl<75> / cell_PIM2
XI19672 bl<31> cbl<15> in1<77> in2<77> sl<31> vdd vss wl<77> / cell_PIM2
XI19671 bl<31> cbl<15> in1<78> in2<78> sl<31> vdd vss wl<78> / cell_PIM2
XI19670 bl<31> cbl<15> in1<79> in2<79> sl<31> vdd vss wl<79> / cell_PIM2
XI19673 bl<31> cbl<15> in1<76> in2<76> sl<31> vdd vss wl<76> / cell_PIM2
XI20843 bl<21> cbl<10> in1<2> in2<2> sl<21> vdd vss wl<2> / cell_PIM2
XI20842 bl<21> cbl<10> in1<1> in2<1> sl<21> vdd vss wl<1> / cell_PIM2
XI19664 bl<29> cbl<14> in1<76> in2<76> sl<29> vdd vss wl<76> / cell_PIM2
XI20208 bl<29> cbl<14> in1<43> in2<43> sl<29> vdd vss wl<43> / cell_PIM2
XI20207 bl<29> cbl<14> in1<42> in2<42> sl<29> vdd vss wl<42> / cell_PIM2
XI20206 bl<29> cbl<14> in1<41> in2<41> sl<29> vdd vss wl<41> / cell_PIM2
XI20205 bl<29> cbl<14> in1<45> in2<45> sl<29> vdd vss wl<45> / cell_PIM2
XI20838 bl<19> cbl<9> in1<0> in2<0> sl<19> vdd vss wl<0> / cell_PIM2
XI20837 bl<19> cbl<9> in1<1> in2<1> sl<19> vdd vss wl<1> / cell_PIM2
XI20836 bl<19> cbl<9> in1<2> in2<2> sl<19> vdd vss wl<2> / cell_PIM2
XI19662 bl<29> cbl<14> in1<79> in2<79> sl<29> vdd vss wl<79> / cell_PIM2
XI19661 bl<29> cbl<14> in1<78> in2<78> sl<29> vdd vss wl<78> / cell_PIM2
XI19660 bl<29> cbl<14> in1<77> in2<77> sl<29> vdd vss wl<77> / cell_PIM2
XI19663 bl<29> cbl<14> in1<75> in2<75> sl<29> vdd vss wl<75> / cell_PIM2
XI20204 bl<29> cbl<14> in1<44> in2<44> sl<29> vdd vss wl<44> / cell_PIM2
XI20832 bl<17> cbl<8> in1<0> in2<0> sl<17> vdd vss wl<0> / cell_PIM2
XI20831 bl<17> cbl<8> in1<2> in2<2> sl<17> vdd vss wl<2> / cell_PIM2
XI20830 bl<17> cbl<8> in1<1> in2<1> sl<17> vdd vss wl<1> / cell_PIM2
XI20826 bl<31> cbl<15> in1<4> in2<4> sl<31> vdd vss wl<4> / cell_PIM2
XI20825 bl<31> cbl<15> in1<3> in2<3> sl<31> vdd vss wl<3> / cell_PIM2
XI20824 bl<31> cbl<15> in1<5> in2<5> sl<31> vdd vss wl<5> / cell_PIM2
XI20198 bl<27> cbl<13> in1<41> in2<41> sl<27> vdd vss wl<41> / cell_PIM2
XI20197 bl<27> cbl<13> in1<42> in2<42> sl<27> vdd vss wl<42> / cell_PIM2
XI19654 bl<27> cbl<13> in1<75> in2<75> sl<27> vdd vss wl<75> / cell_PIM2
XI19652 bl<27> cbl<13> in1<77> in2<77> sl<27> vdd vss wl<77> / cell_PIM2
XI19651 bl<27> cbl<13> in1<78> in2<78> sl<27> vdd vss wl<78> / cell_PIM2
XI19650 bl<27> cbl<13> in1<79> in2<79> sl<27> vdd vss wl<79> / cell_PIM2
XI19653 bl<27> cbl<13> in1<76> in2<76> sl<27> vdd vss wl<76> / cell_PIM2
XI20196 bl<27> cbl<13> in1<43> in2<43> sl<27> vdd vss wl<43> / cell_PIM2
XI20195 bl<27> cbl<13> in1<44> in2<44> sl<27> vdd vss wl<44> / cell_PIM2
XI20194 bl<27> cbl<13> in1<45> in2<45> sl<27> vdd vss wl<45> / cell_PIM2
XI20823 bl<31> cbl<15> in1<6> in2<6> sl<31> vdd vss wl<6> / cell_PIM2
XI20822 bl<31> cbl<15> in1<7> in2<7> sl<31> vdd vss wl<7> / cell_PIM2
XI19644 bl<25> cbl<12> in1<75> in2<75> sl<25> vdd vss wl<75> / cell_PIM2
XI20816 bl<29> cbl<14> in1<3> in2<3> sl<29> vdd vss wl<3> / cell_PIM2
XI20815 bl<29> cbl<14> in1<4> in2<4> sl<29> vdd vss wl<4> / cell_PIM2
XI20814 bl<29> cbl<14> in1<7> in2<7> sl<29> vdd vss wl<7> / cell_PIM2
XI19642 bl<25> cbl<12> in1<77> in2<77> sl<25> vdd vss wl<77> / cell_PIM2
XI19641 bl<25> cbl<12> in1<78> in2<78> sl<25> vdd vss wl<78> / cell_PIM2
XI19640 bl<25> cbl<12> in1<79> in2<79> sl<25> vdd vss wl<79> / cell_PIM2
XI19643 bl<25> cbl<12> in1<76> in2<76> sl<25> vdd vss wl<76> / cell_PIM2
XI20188 bl<25> cbl<12> in1<41> in2<41> sl<25> vdd vss wl<41> / cell_PIM2
XI20187 bl<25> cbl<12> in1<42> in2<42> sl<25> vdd vss wl<42> / cell_PIM2
XI20186 bl<25> cbl<12> in1<43> in2<43> sl<25> vdd vss wl<43> / cell_PIM2
XI20185 bl<25> cbl<12> in1<44> in2<44> sl<25> vdd vss wl<44> / cell_PIM2
XI20813 bl<29> cbl<14> in1<6> in2<6> sl<29> vdd vss wl<6> / cell_PIM2
XI20812 bl<29> cbl<14> in1<5> in2<5> sl<29> vdd vss wl<5> / cell_PIM2
XI20806 bl<27> cbl<13> in1<4> in2<4> sl<27> vdd vss wl<4> / cell_PIM2
XI20805 bl<27> cbl<13> in1<3> in2<3> sl<27> vdd vss wl<3> / cell_PIM2
XI20804 bl<27> cbl<13> in1<5> in2<5> sl<27> vdd vss wl<5> / cell_PIM2
XI20184 bl<25> cbl<12> in1<45> in2<45> sl<25> vdd vss wl<45> / cell_PIM2
XI19634 bl<23> cbl<11> in1<75> in2<75> sl<23> vdd vss wl<75> / cell_PIM2
XI19632 bl<23> cbl<11> in1<77> in2<77> sl<23> vdd vss wl<77> / cell_PIM2
XI19631 bl<23> cbl<11> in1<78> in2<78> sl<23> vdd vss wl<78> / cell_PIM2
XI19630 bl<23> cbl<11> in1<79> in2<79> sl<23> vdd vss wl<79> / cell_PIM2
XI19633 bl<23> cbl<11> in1<76> in2<76> sl<23> vdd vss wl<76> / cell_PIM2
XI20178 bl<23> cbl<11> in1<41> in2<41> sl<23> vdd vss wl<41> / cell_PIM2
XI20177 bl<23> cbl<11> in1<42> in2<42> sl<23> vdd vss wl<42> / cell_PIM2
XI20803 bl<27> cbl<13> in1<6> in2<6> sl<27> vdd vss wl<6> / cell_PIM2
XI20802 bl<27> cbl<13> in1<7> in2<7> sl<27> vdd vss wl<7> / cell_PIM2
XI19624 bl<21> cbl<10> in1<76> in2<76> sl<21> vdd vss wl<76> / cell_PIM2
XI20176 bl<23> cbl<11> in1<43> in2<43> sl<23> vdd vss wl<43> / cell_PIM2
XI20175 bl<23> cbl<11> in1<44> in2<44> sl<23> vdd vss wl<44> / cell_PIM2
XI20174 bl<23> cbl<11> in1<45> in2<45> sl<23> vdd vss wl<45> / cell_PIM2
XI20796 bl<25> cbl<12> in1<4> in2<4> sl<25> vdd vss wl<4> / cell_PIM2
XI20795 bl<25> cbl<12> in1<3> in2<3> sl<25> vdd vss wl<3> / cell_PIM2
XI20794 bl<25> cbl<12> in1<5> in2<5> sl<25> vdd vss wl<5> / cell_PIM2
XI19622 bl<21> cbl<10> in1<79> in2<79> sl<21> vdd vss wl<79> / cell_PIM2
XI19621 bl<21> cbl<10> in1<78> in2<78> sl<21> vdd vss wl<78> / cell_PIM2
XI19620 bl<21> cbl<10> in1<77> in2<77> sl<21> vdd vss wl<77> / cell_PIM2
XI19623 bl<21> cbl<10> in1<75> in2<75> sl<21> vdd vss wl<75> / cell_PIM2
XI20793 bl<25> cbl<12> in1<6> in2<6> sl<25> vdd vss wl<6> / cell_PIM2
XI20792 bl<25> cbl<12> in1<7> in2<7> sl<25> vdd vss wl<7> / cell_PIM2
XI20786 bl<23> cbl<11> in1<4> in2<4> sl<23> vdd vss wl<4> / cell_PIM2
XI20785 bl<23> cbl<11> in1<3> in2<3> sl<23> vdd vss wl<3> / cell_PIM2
XI20784 bl<23> cbl<11> in1<5> in2<5> sl<23> vdd vss wl<5> / cell_PIM2
XI20168 bl<21> cbl<10> in1<43> in2<43> sl<21> vdd vss wl<43> / cell_PIM2
XI20167 bl<21> cbl<10> in1<42> in2<42> sl<21> vdd vss wl<42> / cell_PIM2
XI20166 bl<21> cbl<10> in1<41> in2<41> sl<21> vdd vss wl<41> / cell_PIM2
XI20165 bl<21> cbl<10> in1<45> in2<45> sl<21> vdd vss wl<45> / cell_PIM2
XI19614 bl<19> cbl<9> in1<75> in2<75> sl<19> vdd vss wl<75> / cell_PIM2
XI19612 bl<19> cbl<9> in1<77> in2<77> sl<19> vdd vss wl<77> / cell_PIM2
XI19611 bl<19> cbl<9> in1<78> in2<78> sl<19> vdd vss wl<78> / cell_PIM2
XI19610 bl<19> cbl<9> in1<79> in2<79> sl<19> vdd vss wl<79> / cell_PIM2
XI19613 bl<19> cbl<9> in1<76> in2<76> sl<19> vdd vss wl<76> / cell_PIM2
XI20164 bl<21> cbl<10> in1<44> in2<44> sl<21> vdd vss wl<44> / cell_PIM2
XI20783 bl<23> cbl<11> in1<6> in2<6> sl<23> vdd vss wl<6> / cell_PIM2
XI20782 bl<23> cbl<11> in1<7> in2<7> sl<23> vdd vss wl<7> / cell_PIM2
XI19604 bl<17> cbl<8> in1<76> in2<76> sl<17> vdd vss wl<76> / cell_PIM2
XI20158 bl<19> cbl<9> in1<41> in2<41> sl<19> vdd vss wl<41> / cell_PIM2
XI20157 bl<19> cbl<9> in1<42> in2<42> sl<19> vdd vss wl<42> / cell_PIM2
XI20776 bl<21> cbl<10> in1<3> in2<3> sl<21> vdd vss wl<3> / cell_PIM2
XI20775 bl<21> cbl<10> in1<4> in2<4> sl<21> vdd vss wl<4> / cell_PIM2
XI20774 bl<21> cbl<10> in1<7> in2<7> sl<21> vdd vss wl<7> / cell_PIM2
XI19602 bl<17> cbl<8> in1<79> in2<79> sl<17> vdd vss wl<79> / cell_PIM2
XI19601 bl<17> cbl<8> in1<78> in2<78> sl<17> vdd vss wl<78> / cell_PIM2
XI19600 bl<17> cbl<8> in1<77> in2<77> sl<17> vdd vss wl<77> / cell_PIM2
XI19603 bl<17> cbl<8> in1<75> in2<75> sl<17> vdd vss wl<75> / cell_PIM2
XI20156 bl<19> cbl<9> in1<43> in2<43> sl<19> vdd vss wl<43> / cell_PIM2
XI20155 bl<19> cbl<9> in1<44> in2<44> sl<19> vdd vss wl<44> / cell_PIM2
XI20154 bl<19> cbl<9> in1<45> in2<45> sl<19> vdd vss wl<45> / cell_PIM2
XI20773 bl<21> cbl<10> in1<6> in2<6> sl<21> vdd vss wl<6> / cell_PIM2
XI20772 bl<21> cbl<10> in1<5> in2<5> sl<21> vdd vss wl<5> / cell_PIM2
XI20766 bl<19> cbl<9> in1<4> in2<4> sl<19> vdd vss wl<4> / cell_PIM2
XI20765 bl<19> cbl<9> in1<3> in2<3> sl<19> vdd vss wl<3> / cell_PIM2
XI20764 bl<19> cbl<9> in1<5> in2<5> sl<19> vdd vss wl<5> / cell_PIM2
XI19594 bl<31> cbl<15> in1<80> in2<80> sl<31> vdd vss wl<80> / cell_PIM2
XI19592 bl<31> cbl<15> in1<82> in2<82> sl<31> vdd vss wl<82> / cell_PIM2
XI19591 bl<31> cbl<15> in1<83> in2<83> sl<31> vdd vss wl<83> / cell_PIM2
XI19593 bl<31> cbl<15> in1<81> in2<81> sl<31> vdd vss wl<81> / cell_PIM2
XI20148 bl<17> cbl<8> in1<43> in2<43> sl<17> vdd vss wl<43> / cell_PIM2
XI20147 bl<17> cbl<8> in1<42> in2<42> sl<17> vdd vss wl<42> / cell_PIM2
XI20146 bl<17> cbl<8> in1<41> in2<41> sl<17> vdd vss wl<41> / cell_PIM2
XI20145 bl<17> cbl<8> in1<45> in2<45> sl<17> vdd vss wl<45> / cell_PIM2
XI20763 bl<19> cbl<9> in1<6> in2<6> sl<19> vdd vss wl<6> / cell_PIM2
XI20762 bl<19> cbl<9> in1<7> in2<7> sl<19> vdd vss wl<7> / cell_PIM2
XI19586 bl<29> cbl<14> in1<81> in2<81> sl<29> vdd vss wl<81> / cell_PIM2
XI19585 bl<29> cbl<14> in1<80> in2<80> sl<29> vdd vss wl<80> / cell_PIM2
XI19584 bl<29> cbl<14> in1<83> in2<83> sl<29> vdd vss wl<83> / cell_PIM2
XI20144 bl<17> cbl<8> in1<44> in2<44> sl<17> vdd vss wl<44> / cell_PIM2
XI20756 bl<17> cbl<8> in1<3> in2<3> sl<17> vdd vss wl<3> / cell_PIM2
XI20755 bl<17> cbl<8> in1<4> in2<4> sl<17> vdd vss wl<4> / cell_PIM2
XI20754 bl<17> cbl<8> in1<7> in2<7> sl<17> vdd vss wl<7> / cell_PIM2
XI19583 bl<29> cbl<14> in1<82> in2<82> sl<29> vdd vss wl<82> / cell_PIM2
XI20138 bl<31> cbl<15> in1<46> in2<46> sl<31> vdd vss wl<46> / cell_PIM2
XI20137 bl<31> cbl<15> in1<47> in2<47> sl<31> vdd vss wl<47> / cell_PIM2
XI20753 bl<17> cbl<8> in1<6> in2<6> sl<17> vdd vss wl<6> / cell_PIM2
XI20752 bl<17> cbl<8> in1<5> in2<5> sl<17> vdd vss wl<5> / cell_PIM2
XI20746 bl<31> cbl<15> in1<8> in2<8> sl<31> vdd vss wl<8> / cell_PIM2
XI20745 bl<31> cbl<15> in1<9> in2<9> sl<31> vdd vss wl<9> / cell_PIM2
XI20744 bl<31> cbl<15> in1<10> in2<10> sl<31> vdd vss wl<10> / cell_PIM2
XI20136 bl<31> cbl<15> in1<48> in2<48> sl<31> vdd vss wl<48> / cell_PIM2
XI20135 bl<31> cbl<15> in1<49> in2<49> sl<31> vdd vss wl<49> / cell_PIM2
XI20134 bl<31> cbl<15> in1<50> in2<50> sl<31> vdd vss wl<50> / cell_PIM2
XI19578 bl<27> cbl<13> in1<80> in2<80> sl<27> vdd vss wl<80> / cell_PIM2
XI19577 bl<27> cbl<13> in1<81> in2<81> sl<27> vdd vss wl<81> / cell_PIM2
XI19576 bl<27> cbl<13> in1<82> in2<82> sl<27> vdd vss wl<82> / cell_PIM2
XI19575 bl<27> cbl<13> in1<83> in2<83> sl<27> vdd vss wl<83> / cell_PIM2
XI19570 bl<25> cbl<12> in1<80> in2<80> sl<25> vdd vss wl<80> / cell_PIM2
XI19569 bl<25> cbl<12> in1<81> in2<81> sl<25> vdd vss wl<81> / cell_PIM2
XI20743 bl<31> cbl<15> in1<11> in2<11> sl<31> vdd vss wl<11> / cell_PIM2
XI20742 bl<31> cbl<15> in1<12> in2<12> sl<31> vdd vss wl<12> / cell_PIM2
XI19567 bl<25> cbl<12> in1<83> in2<83> sl<25> vdd vss wl<83> / cell_PIM2
XI19568 bl<25> cbl<12> in1<82> in2<82> sl<25> vdd vss wl<82> / cell_PIM2
XI20128 bl<29> cbl<14> in1<47> in2<47> sl<29> vdd vss wl<47> / cell_PIM2
XI20127 bl<29> cbl<14> in1<46> in2<46> sl<29> vdd vss wl<46> / cell_PIM2
XI20126 bl<29> cbl<14> in1<50> in2<50> sl<29> vdd vss wl<50> / cell_PIM2
XI20125 bl<29> cbl<14> in1<49> in2<49> sl<29> vdd vss wl<49> / cell_PIM2
XI20736 bl<29> cbl<14> in1<9> in2<9> sl<29> vdd vss wl<9> / cell_PIM2
XI20735 bl<29> cbl<14> in1<8> in2<8> sl<29> vdd vss wl<8> / cell_PIM2
XI20734 bl<29> cbl<14> in1<12> in2<12> sl<29> vdd vss wl<12> / cell_PIM2
XI19562 bl<23> cbl<11> in1<80> in2<80> sl<23> vdd vss wl<80> / cell_PIM2
XI19561 bl<23> cbl<11> in1<81> in2<81> sl<23> vdd vss wl<81> / cell_PIM2
XI19560 bl<23> cbl<11> in1<82> in2<82> sl<23> vdd vss wl<82> / cell_PIM2
XI19559 bl<23> cbl<11> in1<83> in2<83> sl<23> vdd vss wl<83> / cell_PIM2
XI20124 bl<29> cbl<14> in1<48> in2<48> sl<29> vdd vss wl<48> / cell_PIM2
XI20733 bl<29> cbl<14> in1<11> in2<11> sl<29> vdd vss wl<11> / cell_PIM2
XI20732 bl<29> cbl<14> in1<10> in2<10> sl<29> vdd vss wl<10> / cell_PIM2
XI20726 bl<27> cbl<13> in1<8> in2<8> sl<27> vdd vss wl<8> / cell_PIM2
XI20725 bl<27> cbl<13> in1<9> in2<9> sl<27> vdd vss wl<9> / cell_PIM2
XI20724 bl<27> cbl<13> in1<10> in2<10> sl<27> vdd vss wl<10> / cell_PIM2
XI20118 bl<27> cbl<13> in1<46> in2<46> sl<27> vdd vss wl<46> / cell_PIM2
XI20117 bl<27> cbl<13> in1<47> in2<47> sl<27> vdd vss wl<47> / cell_PIM2
XI19554 bl<21> cbl<10> in1<81> in2<81> sl<21> vdd vss wl<81> / cell_PIM2
XI19552 bl<21> cbl<10> in1<83> in2<83> sl<21> vdd vss wl<83> / cell_PIM2
XI19551 bl<21> cbl<10> in1<82> in2<82> sl<21> vdd vss wl<82> / cell_PIM2
XI19553 bl<21> cbl<10> in1<80> in2<80> sl<21> vdd vss wl<80> / cell_PIM2
XI20116 bl<27> cbl<13> in1<48> in2<48> sl<27> vdd vss wl<48> / cell_PIM2
XI20115 bl<27> cbl<13> in1<49> in2<49> sl<27> vdd vss wl<49> / cell_PIM2
XI20114 bl<27> cbl<13> in1<50> in2<50> sl<27> vdd vss wl<50> / cell_PIM2
XI20723 bl<27> cbl<13> in1<11> in2<11> sl<27> vdd vss wl<11> / cell_PIM2
XI20722 bl<27> cbl<13> in1<12> in2<12> sl<27> vdd vss wl<12> / cell_PIM2
XI19546 bl<19> cbl<9> in1<80> in2<80> sl<19> vdd vss wl<80> / cell_PIM2
XI19545 bl<19> cbl<9> in1<81> in2<81> sl<19> vdd vss wl<81> / cell_PIM2
XI19544 bl<19> cbl<9> in1<82> in2<82> sl<19> vdd vss wl<82> / cell_PIM2
XI20716 bl<25> cbl<12> in1<8> in2<8> sl<25> vdd vss wl<8> / cell_PIM2
XI20715 bl<25> cbl<12> in1<9> in2<9> sl<25> vdd vss wl<9> / cell_PIM2
XI20714 bl<25> cbl<12> in1<10> in2<10> sl<25> vdd vss wl<10> / cell_PIM2
XI19543 bl<19> cbl<9> in1<83> in2<83> sl<19> vdd vss wl<83> / cell_PIM2
XI20108 bl<25> cbl<12> in1<46> in2<46> sl<25> vdd vss wl<46> / cell_PIM2
XI20107 bl<25> cbl<12> in1<47> in2<47> sl<25> vdd vss wl<47> / cell_PIM2
XI20106 bl<25> cbl<12> in1<48> in2<48> sl<25> vdd vss wl<48> / cell_PIM2
XI20105 bl<25> cbl<12> in1<49> in2<49> sl<25> vdd vss wl<49> / cell_PIM2
XI20713 bl<25> cbl<12> in1<11> in2<11> sl<25> vdd vss wl<11> / cell_PIM2
XI20712 bl<25> cbl<12> in1<12> in2<12> sl<25> vdd vss wl<12> / cell_PIM2
XI20706 bl<23> cbl<11> in1<8> in2<8> sl<23> vdd vss wl<8> / cell_PIM2
XI20705 bl<23> cbl<11> in1<9> in2<9> sl<23> vdd vss wl<9> / cell_PIM2
XI20704 bl<23> cbl<11> in1<10> in2<10> sl<23> vdd vss wl<10> / cell_PIM2
XI20104 bl<25> cbl<12> in1<50> in2<50> sl<25> vdd vss wl<50> / cell_PIM2
XI19538 bl<17> cbl<8> in1<81> in2<81> sl<17> vdd vss wl<81> / cell_PIM2
XI19537 bl<17> cbl<8> in1<80> in2<80> sl<17> vdd vss wl<80> / cell_PIM2
XI19536 bl<17> cbl<8> in1<83> in2<83> sl<17> vdd vss wl<83> / cell_PIM2
XI19535 bl<17> cbl<8> in1<82> in2<82> sl<17> vdd vss wl<82> / cell_PIM2
XI19530 bl<31> cbl<15> in1<84> in2<84> sl<31> vdd vss wl<84> / cell_PIM2
XI19529 bl<31> cbl<15> in1<85> in2<85> sl<31> vdd vss wl<85> / cell_PIM2
XI20098 bl<23> cbl<11> in1<46> in2<46> sl<23> vdd vss wl<46> / cell_PIM2
XI20097 bl<23> cbl<11> in1<47> in2<47> sl<23> vdd vss wl<47> / cell_PIM2
XI20703 bl<23> cbl<11> in1<11> in2<11> sl<23> vdd vss wl<11> / cell_PIM2
XI20702 bl<23> cbl<11> in1<12> in2<12> sl<23> vdd vss wl<12> / cell_PIM2
XI19527 bl<31> cbl<15> in1<87> in2<87> sl<31> vdd vss wl<87> / cell_PIM2
XI19526 bl<31> cbl<15> in1<88> in2<88> sl<31> vdd vss wl<88> / cell_PIM2
XI19528 bl<31> cbl<15> in1<86> in2<86> sl<31> vdd vss wl<86> / cell_PIM2
XI20096 bl<23> cbl<11> in1<48> in2<48> sl<23> vdd vss wl<48> / cell_PIM2
XI20095 bl<23> cbl<11> in1<49> in2<49> sl<23> vdd vss wl<49> / cell_PIM2
XI20094 bl<23> cbl<11> in1<50> in2<50> sl<23> vdd vss wl<50> / cell_PIM2
XI20696 bl<21> cbl<10> in1<9> in2<9> sl<21> vdd vss wl<9> / cell_PIM2
XI20695 bl<21> cbl<10> in1<8> in2<8> sl<21> vdd vss wl<8> / cell_PIM2
XI20694 bl<21> cbl<10> in1<12> in2<12> sl<21> vdd vss wl<12> / cell_PIM2
XI19520 bl<29> cbl<14> in1<86> in2<86> sl<29> vdd vss wl<86> / cell_PIM2
XI19519 bl<29> cbl<14> in1<85> in2<85> sl<29> vdd vss wl<85> / cell_PIM2
XI20693 bl<21> cbl<10> in1<11> in2<11> sl<21> vdd vss wl<11> / cell_PIM2
XI20692 bl<21> cbl<10> in1<10> in2<10> sl<21> vdd vss wl<10> / cell_PIM2
XI20686 bl<19> cbl<9> in1<8> in2<8> sl<19> vdd vss wl<8> / cell_PIM2
XI20685 bl<19> cbl<9> in1<9> in2<9> sl<19> vdd vss wl<9> / cell_PIM2
XI20684 bl<19> cbl<9> in1<10> in2<10> sl<19> vdd vss wl<10> / cell_PIM2
XI20088 bl<21> cbl<10> in1<47> in2<47> sl<21> vdd vss wl<47> / cell_PIM2
XI20087 bl<21> cbl<10> in1<46> in2<46> sl<21> vdd vss wl<46> / cell_PIM2
XI20086 bl<21> cbl<10> in1<50> in2<50> sl<21> vdd vss wl<50> / cell_PIM2
XI20085 bl<21> cbl<10> in1<49> in2<49> sl<21> vdd vss wl<49> / cell_PIM2
XI19518 bl<29> cbl<14> in1<84> in2<84> sl<29> vdd vss wl<84> / cell_PIM2
XI19517 bl<29> cbl<14> in1<88> in2<88> sl<29> vdd vss wl<88> / cell_PIM2
XI19516 bl<29> cbl<14> in1<87> in2<87> sl<29> vdd vss wl<87> / cell_PIM2
XI19510 bl<27> cbl<13> in1<84> in2<84> sl<27> vdd vss wl<84> / cell_PIM2
XI19509 bl<27> cbl<13> in1<85> in2<85> sl<27> vdd vss wl<85> / cell_PIM2
XI20084 bl<21> cbl<10> in1<48> in2<48> sl<21> vdd vss wl<48> / cell_PIM2
XI20683 bl<19> cbl<9> in1<11> in2<11> sl<19> vdd vss wl<11> / cell_PIM2
XI20682 bl<19> cbl<9> in1<12> in2<12> sl<19> vdd vss wl<12> / cell_PIM2
XI19507 bl<27> cbl<13> in1<87> in2<87> sl<27> vdd vss wl<87> / cell_PIM2
XI19506 bl<27> cbl<13> in1<88> in2<88> sl<27> vdd vss wl<88> / cell_PIM2
XI19508 bl<27> cbl<13> in1<86> in2<86> sl<27> vdd vss wl<86> / cell_PIM2
XI20078 bl<19> cbl<9> in1<46> in2<46> sl<19> vdd vss wl<46> / cell_PIM2
XI20077 bl<19> cbl<9> in1<47> in2<47> sl<19> vdd vss wl<47> / cell_PIM2
XI20676 bl<17> cbl<8> in1<9> in2<9> sl<17> vdd vss wl<9> / cell_PIM2
XI20675 bl<17> cbl<8> in1<8> in2<8> sl<17> vdd vss wl<8> / cell_PIM2
XI20674 bl<17> cbl<8> in1<12> in2<12> sl<17> vdd vss wl<12> / cell_PIM2
XI19500 bl<25> cbl<12> in1<84> in2<84> sl<25> vdd vss wl<84> / cell_PIM2
XI19499 bl<25> cbl<12> in1<85> in2<85> sl<25> vdd vss wl<85> / cell_PIM2
XI20076 bl<19> cbl<9> in1<48> in2<48> sl<19> vdd vss wl<48> / cell_PIM2
XI20075 bl<19> cbl<9> in1<49> in2<49> sl<19> vdd vss wl<49> / cell_PIM2
XI20074 bl<19> cbl<9> in1<50> in2<50> sl<19> vdd vss wl<50> / cell_PIM2
XI20673 bl<17> cbl<8> in1<11> in2<11> sl<17> vdd vss wl<11> / cell_PIM2
XI20672 bl<17> cbl<8> in1<10> in2<10> sl<17> vdd vss wl<10> / cell_PIM2
XI20666 bl<31> cbl<15> in1<13> in2<13> sl<31> vdd vss wl<13> / cell_PIM2
XI20665 bl<31> cbl<15> in1<14> in2<14> sl<31> vdd vss wl<14> / cell_PIM2
XI20664 bl<31> cbl<15> in1<15> in2<15> sl<31> vdd vss wl<15> / cell_PIM2
XI19498 bl<25> cbl<12> in1<86> in2<86> sl<25> vdd vss wl<86> / cell_PIM2
XI19497 bl<25> cbl<12> in1<87> in2<87> sl<25> vdd vss wl<87> / cell_PIM2
XI19496 bl<25> cbl<12> in1<88> in2<88> sl<25> vdd vss wl<88> / cell_PIM2
XI19490 bl<23> cbl<11> in1<84> in2<84> sl<23> vdd vss wl<84> / cell_PIM2
XI19489 bl<23> cbl<11> in1<85> in2<85> sl<23> vdd vss wl<85> / cell_PIM2
XI20068 bl<17> cbl<8> in1<47> in2<47> sl<17> vdd vss wl<47> / cell_PIM2
XI20067 bl<17> cbl<8> in1<46> in2<46> sl<17> vdd vss wl<46> / cell_PIM2
XI20066 bl<17> cbl<8> in1<50> in2<50> sl<17> vdd vss wl<50> / cell_PIM2
XI20065 bl<17> cbl<8> in1<49> in2<49> sl<17> vdd vss wl<49> / cell_PIM2
XI20663 bl<31> cbl<15> in1<16> in2<16> sl<31> vdd vss wl<16> / cell_PIM2
XI20662 bl<31> cbl<15> in1<17> in2<17> sl<31> vdd vss wl<17> / cell_PIM2
XI19487 bl<23> cbl<11> in1<87> in2<87> sl<23> vdd vss wl<87> / cell_PIM2
XI19486 bl<23> cbl<11> in1<88> in2<88> sl<23> vdd vss wl<88> / cell_PIM2
XI19488 bl<23> cbl<11> in1<86> in2<86> sl<23> vdd vss wl<86> / cell_PIM2
XI20064 bl<17> cbl<8> in1<48> in2<48> sl<17> vdd vss wl<48> / cell_PIM2
XI20656 bl<29> cbl<14> in1<14> in2<14> sl<29> vdd vss wl<14> / cell_PIM2
XI20655 bl<29> cbl<14> in1<13> in2<13> sl<29> vdd vss wl<13> / cell_PIM2
XI20654 bl<29> cbl<14> in1<17> in2<17> sl<29> vdd vss wl<17> / cell_PIM2
XI19480 bl<21> cbl<10> in1<86> in2<86> sl<21> vdd vss wl<86> / cell_PIM2
XI19479 bl<21> cbl<10> in1<85> in2<85> sl<21> vdd vss wl<85> / cell_PIM2
XI20058 bl<31> cbl<15> in1<51> in2<51> sl<31> vdd vss wl<51> / cell_PIM2
XI20057 bl<31> cbl<15> in1<52> in2<52> sl<31> vdd vss wl<52> / cell_PIM2
XI20653 bl<29> cbl<14> in1<16> in2<16> sl<29> vdd vss wl<16> / cell_PIM2
XI20652 bl<29> cbl<14> in1<15> in2<15> sl<29> vdd vss wl<15> / cell_PIM2
XI20646 bl<27> cbl<13> in1<13> in2<13> sl<27> vdd vss wl<13> / cell_PIM2
XI20645 bl<27> cbl<13> in1<14> in2<14> sl<27> vdd vss wl<14> / cell_PIM2
XI20644 bl<27> cbl<13> in1<15> in2<15> sl<27> vdd vss wl<15> / cell_PIM2
XI20056 bl<31> cbl<15> in1<53> in2<53> sl<31> vdd vss wl<53> / cell_PIM2
XI20055 bl<31> cbl<15> in1<54> in2<54> sl<31> vdd vss wl<54> / cell_PIM2
XI20054 bl<31> cbl<15> in1<55> in2<55> sl<31> vdd vss wl<55> / cell_PIM2
XI19478 bl<21> cbl<10> in1<84> in2<84> sl<21> vdd vss wl<84> / cell_PIM2
XI19477 bl<21> cbl<10> in1<88> in2<88> sl<21> vdd vss wl<88> / cell_PIM2
XI19476 bl<21> cbl<10> in1<87> in2<87> sl<21> vdd vss wl<87> / cell_PIM2
XI19470 bl<19> cbl<9> in1<84> in2<84> sl<19> vdd vss wl<84> / cell_PIM2
XI19469 bl<19> cbl<9> in1<85> in2<85> sl<19> vdd vss wl<85> / cell_PIM2
XI20643 bl<27> cbl<13> in1<16> in2<16> sl<27> vdd vss wl<16> / cell_PIM2
XI20642 bl<27> cbl<13> in1<17> in2<17> sl<27> vdd vss wl<17> / cell_PIM2
XI19467 bl<19> cbl<9> in1<87> in2<87> sl<19> vdd vss wl<87> / cell_PIM2
XI19466 bl<19> cbl<9> in1<88> in2<88> sl<19> vdd vss wl<88> / cell_PIM2
XI19468 bl<19> cbl<9> in1<86> in2<86> sl<19> vdd vss wl<86> / cell_PIM2
XI20048 bl<29> cbl<14> in1<52> in2<52> sl<29> vdd vss wl<52> / cell_PIM2
XI20047 bl<29> cbl<14> in1<51> in2<51> sl<29> vdd vss wl<51> / cell_PIM2
XI20046 bl<29> cbl<14> in1<55> in2<55> sl<29> vdd vss wl<55> / cell_PIM2
XI20045 bl<29> cbl<14> in1<54> in2<54> sl<29> vdd vss wl<54> / cell_PIM2
XI20636 bl<25> cbl<12> in1<13> in2<13> sl<25> vdd vss wl<13> / cell_PIM2
XI20635 bl<25> cbl<12> in1<14> in2<14> sl<25> vdd vss wl<14> / cell_PIM2
XI20634 bl<25> cbl<12> in1<15> in2<15> sl<25> vdd vss wl<15> / cell_PIM2
XI19460 bl<17> cbl<8> in1<86> in2<86> sl<17> vdd vss wl<86> / cell_PIM2
XI19459 bl<17> cbl<8> in1<85> in2<85> sl<17> vdd vss wl<85> / cell_PIM2
XI20044 bl<29> cbl<14> in1<53> in2<53> sl<29> vdd vss wl<53> / cell_PIM2
XI20633 bl<25> cbl<12> in1<16> in2<16> sl<25> vdd vss wl<16> / cell_PIM2
XI20632 bl<25> cbl<12> in1<17> in2<17> sl<25> vdd vss wl<17> / cell_PIM2
XI20626 bl<23> cbl<11> in1<13> in2<13> sl<23> vdd vss wl<13> / cell_PIM2
XI20625 bl<23> cbl<11> in1<14> in2<14> sl<23> vdd vss wl<14> / cell_PIM2
XI20624 bl<23> cbl<11> in1<15> in2<15> sl<23> vdd vss wl<15> / cell_PIM2
XI20038 bl<27> cbl<13> in1<51> in2<51> sl<27> vdd vss wl<51> / cell_PIM2
XI20037 bl<27> cbl<13> in1<52> in2<52> sl<27> vdd vss wl<52> / cell_PIM2
XI19458 bl<17> cbl<8> in1<84> in2<84> sl<17> vdd vss wl<84> / cell_PIM2
XI19457 bl<17> cbl<8> in1<88> in2<88> sl<17> vdd vss wl<88> / cell_PIM2
XI19456 bl<17> cbl<8> in1<87> in2<87> sl<17> vdd vss wl<87> / cell_PIM2
XI19450 bl<31> cbl<15> in1<89> in2<89> sl<31> vdd vss wl<89> / cell_PIM2
XI19449 bl<31> cbl<15> in1<90> in2<90> sl<31> vdd vss wl<90> / cell_PIM2
XI20036 bl<27> cbl<13> in1<53> in2<53> sl<27> vdd vss wl<53> / cell_PIM2
XI20035 bl<27> cbl<13> in1<54> in2<54> sl<27> vdd vss wl<54> / cell_PIM2
XI20034 bl<27> cbl<13> in1<55> in2<55> sl<27> vdd vss wl<55> / cell_PIM2
XI20623 bl<23> cbl<11> in1<16> in2<16> sl<23> vdd vss wl<16> / cell_PIM2
XI20622 bl<23> cbl<11> in1<17> in2<17> sl<23> vdd vss wl<17> / cell_PIM2
XI19447 bl<31> cbl<15> in1<92> in2<92> sl<31> vdd vss wl<92> / cell_PIM2
XI19446 bl<31> cbl<15> in1<93> in2<93> sl<31> vdd vss wl<93> / cell_PIM2
XI19448 bl<31> cbl<15> in1<91> in2<91> sl<31> vdd vss wl<91> / cell_PIM2
XI20616 bl<21> cbl<10> in1<14> in2<14> sl<21> vdd vss wl<14> / cell_PIM2
XI20615 bl<21> cbl<10> in1<13> in2<13> sl<21> vdd vss wl<13> / cell_PIM2
XI20614 bl<21> cbl<10> in1<17> in2<17> sl<21> vdd vss wl<17> / cell_PIM2
XI17813 bl<11> cbl<5> in1<126> in2<126> sl<11> vdd vss wl<126> / cell_PIM2
XI17812 bl<11> cbl<5> in1<125> in2<125> sl<11> vdd vss wl<125> / cell_PIM2
XI18463 bl<13> cbl<6> in1<44> in2<44> sl<13> vdd vss wl<44> / cell_PIM2
XI19113 bl<25> cbl<12> in1<111> in2<111> sl<25> vdd vss wl<111> / cell_PIM2
XI19112 bl<25> cbl<12> in1<112> in2<112> sl<25> vdd vss wl<112> / cell_PIM2
XI19106 bl<23> cbl<11> in1<108> in2<108> sl<23> vdd vss wl<108> / cell_PIM2
XI19105 bl<23> cbl<11> in1<109> in2<109> sl<23> vdd vss wl<109> / cell_PIM2
XI19104 bl<23> cbl<11> in1<110> in2<110> sl<23> vdd vss wl<110> / cell_PIM2
XI18458 bl<11> cbl<5> in1<44> in2<44> sl<11> vdd vss wl<44> / cell_PIM2
XI18457 bl<11> cbl<5> in1<45> in2<45> sl<11> vdd vss wl<45> / cell_PIM2
XI18456 bl<11> cbl<5> in1<46> in2<46> sl<11> vdd vss wl<46> / cell_PIM2
XI18455 bl<11> cbl<5> in1<47> in2<47> sl<11> vdd vss wl<47> / cell_PIM2
XI17808 bl<9> cbl<4> in1<127> in2<127> sl<9> vdd vss wl<127> / cell_PIM2
XI17807 bl<9> cbl<4> in1<126> in2<126> sl<9> vdd vss wl<126> / cell_PIM2
XI17806 bl<9> cbl<4> in1<125> in2<125> sl<9> vdd vss wl<125> / cell_PIM2
XI17802 bl<7> cbl<3> in1<0> in2<0> sl<7> vdd vss wl<0> / cell_PIM2
XI17800 bl<5> cbl<2> in1<0> in2<0> sl<5> vdd vss wl<0> / cell_PIM2
XI18450 bl<9> cbl<4> in1<47> in2<47> sl<9> vdd vss wl<47> / cell_PIM2
XI18449 bl<9> cbl<4> in1<46> in2<46> sl<9> vdd vss wl<46> / cell_PIM2
XI19103 bl<23> cbl<11> in1<111> in2<111> sl<23> vdd vss wl<111> / cell_PIM2
XI19102 bl<23> cbl<11> in1<112> in2<112> sl<23> vdd vss wl<112> / cell_PIM2
XI17798 bl<7> cbl<3> in1<1> in2<1> sl<7> vdd vss wl<1> / cell_PIM2
XI17797 bl<7> cbl<3> in1<4> in2<4> sl<7> vdd vss wl<4> / cell_PIM2
XI17796 bl<7> cbl<3> in1<3> in2<3> sl<7> vdd vss wl<3> / cell_PIM2
XI17795 bl<7> cbl<3> in1<2> in2<2> sl<7> vdd vss wl<2> / cell_PIM2
XI18448 bl<9> cbl<4> in1<45> in2<45> sl<9> vdd vss wl<45> / cell_PIM2
XI18447 bl<9> cbl<4> in1<44> in2<44> sl<9> vdd vss wl<44> / cell_PIM2
XI19096 bl<21> cbl<10> in1<110> in2<110> sl<21> vdd vss wl<110> / cell_PIM2
XI19095 bl<21> cbl<10> in1<109> in2<109> sl<21> vdd vss wl<109> / cell_PIM2
XI19094 bl<21> cbl<10> in1<108> in2<108> sl<21> vdd vss wl<108> / cell_PIM2
XI17790 bl<5> cbl<2> in1<2> in2<2> sl<5> vdd vss wl<2> / cell_PIM2
XI17789 bl<5> cbl<2> in1<3> in2<3> sl<5> vdd vss wl<3> / cell_PIM2
XI18442 bl<15> cbl<7> in1<48> in2<48> sl<15> vdd vss wl<48> / cell_PIM2
XI18441 bl<15> cbl<7> in1<49> in2<49> sl<15> vdd vss wl<49> / cell_PIM2
XI18440 bl<15> cbl<7> in1<50> in2<50> sl<15> vdd vss wl<50> / cell_PIM2
XI18439 bl<15> cbl<7> in1<51> in2<51> sl<15> vdd vss wl<51> / cell_PIM2
XI19093 bl<21> cbl<10> in1<112> in2<112> sl<21> vdd vss wl<112> / cell_PIM2
XI19092 bl<21> cbl<10> in1<111> in2<111> sl<21> vdd vss wl<111> / cell_PIM2
XI19086 bl<19> cbl<9> in1<108> in2<108> sl<19> vdd vss wl<108> / cell_PIM2
XI19085 bl<19> cbl<9> in1<109> in2<109> sl<19> vdd vss wl<109> / cell_PIM2
XI19084 bl<19> cbl<9> in1<110> in2<110> sl<19> vdd vss wl<110> / cell_PIM2
XI18438 bl<15> cbl<7> in1<52> in2<52> sl<15> vdd vss wl<52> / cell_PIM2
XI17788 bl<5> cbl<2> in1<4> in2<4> sl<5> vdd vss wl<4> / cell_PIM2
XI17787 bl<5> cbl<2> in1<1> in2<1> sl<5> vdd vss wl<1> / cell_PIM2
XI17782 bl<7> cbl<3> in1<5> in2<5> sl<7> vdd vss wl<5> / cell_PIM2
XI17781 bl<7> cbl<3> in1<6> in2<6> sl<7> vdd vss wl<6> / cell_PIM2
XI17780 bl<7> cbl<3> in1<7> in2<7> sl<7> vdd vss wl<7> / cell_PIM2
XI17779 bl<7> cbl<3> in1<8> in2<8> sl<7> vdd vss wl<8> / cell_PIM2
XI18432 bl<13> cbl<6> in1<52> in2<52> sl<13> vdd vss wl<52> / cell_PIM2
XI18431 bl<13> cbl<6> in1<51> in2<51> sl<13> vdd vss wl<51> / cell_PIM2
XI18430 bl<13> cbl<6> in1<50> in2<50> sl<13> vdd vss wl<50> / cell_PIM2
XI18429 bl<13> cbl<6> in1<49> in2<49> sl<13> vdd vss wl<49> / cell_PIM2
XI19083 bl<19> cbl<9> in1<111> in2<111> sl<19> vdd vss wl<111> / cell_PIM2
XI19082 bl<19> cbl<9> in1<112> in2<112> sl<19> vdd vss wl<112> / cell_PIM2
XI17778 bl<7> cbl<3> in1<9> in2<9> sl<7> vdd vss wl<9> / cell_PIM2
XI18428 bl<13> cbl<6> in1<48> in2<48> sl<13> vdd vss wl<48> / cell_PIM2
XI19076 bl<17> cbl<8> in1<110> in2<110> sl<17> vdd vss wl<110> / cell_PIM2
XI19075 bl<17> cbl<8> in1<109> in2<109> sl<17> vdd vss wl<109> / cell_PIM2
XI19074 bl<17> cbl<8> in1<108> in2<108> sl<17> vdd vss wl<108> / cell_PIM2
XI17772 bl<5> cbl<2> in1<9> in2<9> sl<5> vdd vss wl<9> / cell_PIM2
XI17771 bl<5> cbl<2> in1<8> in2<8> sl<5> vdd vss wl<8> / cell_PIM2
XI17770 bl<5> cbl<2> in1<7> in2<7> sl<5> vdd vss wl<7> / cell_PIM2
XI17769 bl<5> cbl<2> in1<6> in2<6> sl<5> vdd vss wl<6> / cell_PIM2
XI18422 bl<11> cbl<5> in1<48> in2<48> sl<11> vdd vss wl<48> / cell_PIM2
XI18421 bl<11> cbl<5> in1<49> in2<49> sl<11> vdd vss wl<49> / cell_PIM2
XI18420 bl<11> cbl<5> in1<50> in2<50> sl<11> vdd vss wl<50> / cell_PIM2
XI18419 bl<11> cbl<5> in1<51> in2<51> sl<11> vdd vss wl<51> / cell_PIM2
XI19073 bl<17> cbl<8> in1<112> in2<112> sl<17> vdd vss wl<112> / cell_PIM2
XI19072 bl<17> cbl<8> in1<111> in2<111> sl<17> vdd vss wl<111> / cell_PIM2
XI19066 bl<31> cbl<15> in1<113> in2<113> sl<31> vdd vss wl<113> / cell_PIM2
XI19065 bl<31> cbl<15> in1<114> in2<114> sl<31> vdd vss wl<114> / cell_PIM2
XI19064 bl<31> cbl<15> in1<115> in2<115> sl<31> vdd vss wl<115> / cell_PIM2
XI18418 bl<11> cbl<5> in1<52> in2<52> sl<11> vdd vss wl<52> / cell_PIM2
XI17768 bl<5> cbl<2> in1<5> in2<5> sl<5> vdd vss wl<5> / cell_PIM2
XI17762 bl<7> cbl<3> in1<10> in2<10> sl<7> vdd vss wl<10> / cell_PIM2
XI17761 bl<7> cbl<3> in1<11> in2<11> sl<7> vdd vss wl<11> / cell_PIM2
XI17760 bl<7> cbl<3> in1<12> in2<12> sl<7> vdd vss wl<12> / cell_PIM2
XI17759 bl<7> cbl<3> in1<13> in2<13> sl<7> vdd vss wl<13> / cell_PIM2
XI18412 bl<9> cbl<4> in1<52> in2<52> sl<9> vdd vss wl<52> / cell_PIM2
XI18411 bl<9> cbl<4> in1<51> in2<51> sl<9> vdd vss wl<51> / cell_PIM2
XI18410 bl<9> cbl<4> in1<50> in2<50> sl<9> vdd vss wl<50> / cell_PIM2
XI18409 bl<9> cbl<4> in1<49> in2<49> sl<9> vdd vss wl<49> / cell_PIM2
XI19063 bl<31> cbl<15> in1<116> in2<116> sl<31> vdd vss wl<116> / cell_PIM2
XI19062 bl<31> cbl<15> in1<117> in2<117> sl<31> vdd vss wl<117> / cell_PIM2
XI17758 bl<7> cbl<3> in1<14> in2<14> sl<7> vdd vss wl<14> / cell_PIM2
XI18408 bl<9> cbl<4> in1<48> in2<48> sl<9> vdd vss wl<48> / cell_PIM2
XI19056 bl<29> cbl<14> in1<115> in2<115> sl<29> vdd vss wl<115> / cell_PIM2
XI19055 bl<29> cbl<14> in1<114> in2<114> sl<29> vdd vss wl<114> / cell_PIM2
XI19054 bl<29> cbl<14> in1<113> in2<113> sl<29> vdd vss wl<113> / cell_PIM2
XI17752 bl<5> cbl<2> in1<14> in2<14> sl<5> vdd vss wl<14> / cell_PIM2
XI17751 bl<5> cbl<2> in1<13> in2<13> sl<5> vdd vss wl<13> / cell_PIM2
XI17750 bl<5> cbl<2> in1<12> in2<12> sl<5> vdd vss wl<12> / cell_PIM2
XI17749 bl<5> cbl<2> in1<11> in2<11> sl<5> vdd vss wl<11> / cell_PIM2
XI18402 bl<15> cbl<7> in1<53> in2<53> sl<15> vdd vss wl<53> / cell_PIM2
XI18401 bl<15> cbl<7> in1<54> in2<54> sl<15> vdd vss wl<54> / cell_PIM2
XI18400 bl<15> cbl<7> in1<55> in2<55> sl<15> vdd vss wl<55> / cell_PIM2
XI18399 bl<15> cbl<7> in1<56> in2<56> sl<15> vdd vss wl<56> / cell_PIM2
XI19053 bl<29> cbl<14> in1<117> in2<117> sl<29> vdd vss wl<117> / cell_PIM2
XI19052 bl<29> cbl<14> in1<116> in2<116> sl<29> vdd vss wl<116> / cell_PIM2
XI19046 bl<27> cbl<13> in1<113> in2<113> sl<27> vdd vss wl<113> / cell_PIM2
XI19045 bl<27> cbl<13> in1<114> in2<114> sl<27> vdd vss wl<114> / cell_PIM2
XI19044 bl<27> cbl<13> in1<115> in2<115> sl<27> vdd vss wl<115> / cell_PIM2
XI18398 bl<15> cbl<7> in1<57> in2<57> sl<15> vdd vss wl<57> / cell_PIM2
XI17748 bl<5> cbl<2> in1<10> in2<10> sl<5> vdd vss wl<10> / cell_PIM2
XI17742 bl<7> cbl<3> in1<15> in2<15> sl<7> vdd vss wl<15> / cell_PIM2
XI17741 bl<7> cbl<3> in1<16> in2<16> sl<7> vdd vss wl<16> / cell_PIM2
XI17740 bl<7> cbl<3> in1<17> in2<17> sl<7> vdd vss wl<17> / cell_PIM2
XI17739 bl<7> cbl<3> in1<18> in2<18> sl<7> vdd vss wl<18> / cell_PIM2
XI18392 bl<13> cbl<6> in1<57> in2<57> sl<13> vdd vss wl<57> / cell_PIM2
XI18391 bl<13> cbl<6> in1<56> in2<56> sl<13> vdd vss wl<56> / cell_PIM2
XI18390 bl<13> cbl<6> in1<55> in2<55> sl<13> vdd vss wl<55> / cell_PIM2
XI18389 bl<13> cbl<6> in1<54> in2<54> sl<13> vdd vss wl<54> / cell_PIM2
XI19043 bl<27> cbl<13> in1<116> in2<116> sl<27> vdd vss wl<116> / cell_PIM2
XI19042 bl<27> cbl<13> in1<117> in2<117> sl<27> vdd vss wl<117> / cell_PIM2
XI17738 bl<7> cbl<3> in1<19> in2<19> sl<7> vdd vss wl<19> / cell_PIM2
XI18388 bl<13> cbl<6> in1<53> in2<53> sl<13> vdd vss wl<53> / cell_PIM2
XI19036 bl<25> cbl<12> in1<113> in2<113> sl<25> vdd vss wl<113> / cell_PIM2
XI19035 bl<25> cbl<12> in1<114> in2<114> sl<25> vdd vss wl<114> / cell_PIM2
XI19034 bl<25> cbl<12> in1<115> in2<115> sl<25> vdd vss wl<115> / cell_PIM2
XI17732 bl<5> cbl<2> in1<19> in2<19> sl<5> vdd vss wl<19> / cell_PIM2
XI17731 bl<5> cbl<2> in1<18> in2<18> sl<5> vdd vss wl<18> / cell_PIM2
XI17730 bl<5> cbl<2> in1<17> in2<17> sl<5> vdd vss wl<17> / cell_PIM2
XI17729 bl<5> cbl<2> in1<16> in2<16> sl<5> vdd vss wl<16> / cell_PIM2
XI18382 bl<11> cbl<5> in1<53> in2<53> sl<11> vdd vss wl<53> / cell_PIM2
XI18381 bl<11> cbl<5> in1<54> in2<54> sl<11> vdd vss wl<54> / cell_PIM2
XI18380 bl<11> cbl<5> in1<55> in2<55> sl<11> vdd vss wl<55> / cell_PIM2
XI18379 bl<11> cbl<5> in1<56> in2<56> sl<11> vdd vss wl<56> / cell_PIM2
XI19033 bl<25> cbl<12> in1<116> in2<116> sl<25> vdd vss wl<116> / cell_PIM2
XI19032 bl<25> cbl<12> in1<117> in2<117> sl<25> vdd vss wl<117> / cell_PIM2
XI19026 bl<23> cbl<11> in1<113> in2<113> sl<23> vdd vss wl<113> / cell_PIM2
XI19025 bl<23> cbl<11> in1<114> in2<114> sl<23> vdd vss wl<114> / cell_PIM2
XI19024 bl<23> cbl<11> in1<115> in2<115> sl<23> vdd vss wl<115> / cell_PIM2
XI18378 bl<11> cbl<5> in1<57> in2<57> sl<11> vdd vss wl<57> / cell_PIM2
XI17728 bl<5> cbl<2> in1<15> in2<15> sl<5> vdd vss wl<15> / cell_PIM2
XI17722 bl<7> cbl<3> in1<20> in2<20> sl<7> vdd vss wl<20> / cell_PIM2
XI17721 bl<7> cbl<3> in1<21> in2<21> sl<7> vdd vss wl<21> / cell_PIM2
XI17720 bl<7> cbl<3> in1<22> in2<22> sl<7> vdd vss wl<22> / cell_PIM2
XI17719 bl<7> cbl<3> in1<23> in2<23> sl<7> vdd vss wl<23> / cell_PIM2
XI18372 bl<9> cbl<4> in1<57> in2<57> sl<9> vdd vss wl<57> / cell_PIM2
XI18371 bl<9> cbl<4> in1<56> in2<56> sl<9> vdd vss wl<56> / cell_PIM2
XI18370 bl<9> cbl<4> in1<55> in2<55> sl<9> vdd vss wl<55> / cell_PIM2
XI18369 bl<9> cbl<4> in1<54> in2<54> sl<9> vdd vss wl<54> / cell_PIM2
XI19023 bl<23> cbl<11> in1<116> in2<116> sl<23> vdd vss wl<116> / cell_PIM2
XI19022 bl<23> cbl<11> in1<117> in2<117> sl<23> vdd vss wl<117> / cell_PIM2
XI17718 bl<7> cbl<3> in1<24> in2<24> sl<7> vdd vss wl<24> / cell_PIM2
XI18368 bl<9> cbl<4> in1<53> in2<53> sl<9> vdd vss wl<53> / cell_PIM2
XI19016 bl<21> cbl<10> in1<115> in2<115> sl<21> vdd vss wl<115> / cell_PIM2
XI19015 bl<21> cbl<10> in1<114> in2<114> sl<21> vdd vss wl<114> / cell_PIM2
XI19014 bl<21> cbl<10> in1<113> in2<113> sl<21> vdd vss wl<113> / cell_PIM2
XI17712 bl<5> cbl<2> in1<24> in2<24> sl<5> vdd vss wl<24> / cell_PIM2
XI17711 bl<5> cbl<2> in1<23> in2<23> sl<5> vdd vss wl<23> / cell_PIM2
XI17710 bl<5> cbl<2> in1<22> in2<22> sl<5> vdd vss wl<22> / cell_PIM2
XI17709 bl<5> cbl<2> in1<21> in2<21> sl<5> vdd vss wl<21> / cell_PIM2
XI18362 bl<15> cbl<7> in1<58> in2<58> sl<15> vdd vss wl<58> / cell_PIM2
XI18361 bl<15> cbl<7> in1<59> in2<59> sl<15> vdd vss wl<59> / cell_PIM2
XI18360 bl<15> cbl<7> in1<60> in2<60> sl<15> vdd vss wl<60> / cell_PIM2
XI18359 bl<15> cbl<7> in1<61> in2<61> sl<15> vdd vss wl<61> / cell_PIM2
XI19013 bl<21> cbl<10> in1<117> in2<117> sl<21> vdd vss wl<117> / cell_PIM2
XI19012 bl<21> cbl<10> in1<116> in2<116> sl<21> vdd vss wl<116> / cell_PIM2
XI19006 bl<19> cbl<9> in1<113> in2<113> sl<19> vdd vss wl<113> / cell_PIM2
XI19005 bl<19> cbl<9> in1<114> in2<114> sl<19> vdd vss wl<114> / cell_PIM2
XI19004 bl<19> cbl<9> in1<115> in2<115> sl<19> vdd vss wl<115> / cell_PIM2
XI18358 bl<15> cbl<7> in1<62> in2<62> sl<15> vdd vss wl<62> / cell_PIM2
XI17708 bl<5> cbl<2> in1<20> in2<20> sl<5> vdd vss wl<20> / cell_PIM2
XI17702 bl<7> cbl<3> in1<25> in2<25> sl<7> vdd vss wl<25> / cell_PIM2
XI17701 bl<7> cbl<3> in1<26> in2<26> sl<7> vdd vss wl<26> / cell_PIM2
XI17700 bl<7> cbl<3> in1<27> in2<27> sl<7> vdd vss wl<27> / cell_PIM2
XI17699 bl<7> cbl<3> in1<28> in2<28> sl<7> vdd vss wl<28> / cell_PIM2
XI18352 bl<13> cbl<6> in1<62> in2<62> sl<13> vdd vss wl<62> / cell_PIM2
XI18351 bl<13> cbl<6> in1<61> in2<61> sl<13> vdd vss wl<61> / cell_PIM2
XI18350 bl<13> cbl<6> in1<60> in2<60> sl<13> vdd vss wl<60> / cell_PIM2
XI18349 bl<13> cbl<6> in1<59> in2<59> sl<13> vdd vss wl<59> / cell_PIM2
XI19003 bl<19> cbl<9> in1<116> in2<116> sl<19> vdd vss wl<116> / cell_PIM2
XI19002 bl<19> cbl<9> in1<117> in2<117> sl<19> vdd vss wl<117> / cell_PIM2
XI17694 bl<5> cbl<2> in1<28> in2<28> sl<5> vdd vss wl<28> / cell_PIM2
XI18348 bl<13> cbl<6> in1<58> in2<58> sl<13> vdd vss wl<58> / cell_PIM2
XI18996 bl<17> cbl<8> in1<115> in2<115> sl<17> vdd vss wl<115> / cell_PIM2
XI18995 bl<17> cbl<8> in1<114> in2<114> sl<17> vdd vss wl<114> / cell_PIM2
XI18994 bl<17> cbl<8> in1<113> in2<113> sl<17> vdd vss wl<113> / cell_PIM2
XI17693 bl<5> cbl<2> in1<27> in2<27> sl<5> vdd vss wl<27> / cell_PIM2
XI17692 bl<5> cbl<2> in1<26> in2<26> sl<5> vdd vss wl<26> / cell_PIM2
XI17691 bl<5> cbl<2> in1<25> in2<25> sl<5> vdd vss wl<25> / cell_PIM2
XI18342 bl<11> cbl<5> in1<58> in2<58> sl<11> vdd vss wl<58> / cell_PIM2
XI18341 bl<11> cbl<5> in1<59> in2<59> sl<11> vdd vss wl<59> / cell_PIM2
XI18340 bl<11> cbl<5> in1<60> in2<60> sl<11> vdd vss wl<60> / cell_PIM2
XI18339 bl<11> cbl<5> in1<61> in2<61> sl<11> vdd vss wl<61> / cell_PIM2
XI18993 bl<17> cbl<8> in1<117> in2<117> sl<17> vdd vss wl<117> / cell_PIM2
XI18992 bl<17> cbl<8> in1<116> in2<116> sl<17> vdd vss wl<116> / cell_PIM2
XI18986 bl<31> cbl<15> in1<118> in2<118> sl<31> vdd vss wl<118> / cell_PIM2
XI18985 bl<31> cbl<15> in1<119> in2<119> sl<31> vdd vss wl<119> / cell_PIM2
XI18984 bl<31> cbl<15> in1<120> in2<120> sl<31> vdd vss wl<120> / cell_PIM2
XI18338 bl<11> cbl<5> in1<62> in2<62> sl<11> vdd vss wl<62> / cell_PIM2
XI17686 bl<7> cbl<3> in1<29> in2<29> sl<7> vdd vss wl<29> / cell_PIM2
XI17685 bl<7> cbl<3> in1<30> in2<30> sl<7> vdd vss wl<30> / cell_PIM2
XI17684 bl<7> cbl<3> in1<31> in2<31> sl<7> vdd vss wl<31> / cell_PIM2
XI17683 bl<7> cbl<3> in1<32> in2<32> sl<7> vdd vss wl<32> / cell_PIM2
XI17682 bl<7> cbl<3> in1<33> in2<33> sl<7> vdd vss wl<33> / cell_PIM2
XI18332 bl<9> cbl<4> in1<62> in2<62> sl<9> vdd vss wl<62> / cell_PIM2
XI18331 bl<9> cbl<4> in1<61> in2<61> sl<9> vdd vss wl<61> / cell_PIM2
XI18330 bl<9> cbl<4> in1<60> in2<60> sl<9> vdd vss wl<60> / cell_PIM2
XI18329 bl<9> cbl<4> in1<59> in2<59> sl<9> vdd vss wl<59> / cell_PIM2
XI18983 bl<31> cbl<15> in1<121> in2<121> sl<31> vdd vss wl<121> / cell_PIM2
XI18982 bl<31> cbl<15> in1<122> in2<122> sl<31> vdd vss wl<122> / cell_PIM2
XI17676 bl<5> cbl<2> in1<33> in2<33> sl<5> vdd vss wl<33> / cell_PIM2
XI17675 bl<5> cbl<2> in1<32> in2<32> sl<5> vdd vss wl<32> / cell_PIM2
XI17674 bl<5> cbl<2> in1<31> in2<31> sl<5> vdd vss wl<31> / cell_PIM2
XI18328 bl<9> cbl<4> in1<58> in2<58> sl<9> vdd vss wl<58> / cell_PIM2
XI18976 bl<29> cbl<14> in1<119> in2<119> sl<29> vdd vss wl<119> / cell_PIM2
XI18975 bl<29> cbl<14> in1<118> in2<118> sl<29> vdd vss wl<118> / cell_PIM2
XI18974 bl<29> cbl<14> in1<122> in2<122> sl<29> vdd vss wl<122> / cell_PIM2
XI17673 bl<5> cbl<2> in1<30> in2<30> sl<5> vdd vss wl<30> / cell_PIM2
XI17672 bl<5> cbl<2> in1<29> in2<29> sl<5> vdd vss wl<29> / cell_PIM2
XI18322 bl<15> cbl<7> in1<63> in2<63> sl<15> vdd vss wl<63> / cell_PIM2
XI18321 bl<15> cbl<7> in1<64> in2<64> sl<15> vdd vss wl<64> / cell_PIM2
XI18320 bl<15> cbl<7> in1<65> in2<65> sl<15> vdd vss wl<65> / cell_PIM2
XI18319 bl<15> cbl<7> in1<66> in2<66> sl<15> vdd vss wl<66> / cell_PIM2
XI18973 bl<29> cbl<14> in1<121> in2<121> sl<29> vdd vss wl<121> / cell_PIM2
XI18972 bl<29> cbl<14> in1<120> in2<120> sl<29> vdd vss wl<120> / cell_PIM2
XI18966 bl<27> cbl<13> in1<118> in2<118> sl<27> vdd vss wl<118> / cell_PIM2
XI18965 bl<27> cbl<13> in1<119> in2<119> sl<27> vdd vss wl<119> / cell_PIM2
XI18964 bl<27> cbl<13> in1<120> in2<120> sl<27> vdd vss wl<120> / cell_PIM2
XI18318 bl<15> cbl<7> in1<67> in2<67> sl<15> vdd vss wl<67> / cell_PIM2
XI17666 bl<7> cbl<3> in1<34> in2<34> sl<7> vdd vss wl<34> / cell_PIM2
XI17665 bl<7> cbl<3> in1<35> in2<35> sl<7> vdd vss wl<35> / cell_PIM2
XI17664 bl<7> cbl<3> in1<36> in2<36> sl<7> vdd vss wl<36> / cell_PIM2
XI17663 bl<7> cbl<3> in1<37> in2<37> sl<7> vdd vss wl<37> / cell_PIM2
XI17662 bl<7> cbl<3> in1<38> in2<38> sl<7> vdd vss wl<38> / cell_PIM2
XI18312 bl<13> cbl<6> in1<67> in2<67> sl<13> vdd vss wl<67> / cell_PIM2
XI18311 bl<13> cbl<6> in1<66> in2<66> sl<13> vdd vss wl<66> / cell_PIM2
XI18310 bl<13> cbl<6> in1<65> in2<65> sl<13> vdd vss wl<65> / cell_PIM2
XI18309 bl<13> cbl<6> in1<64> in2<64> sl<13> vdd vss wl<64> / cell_PIM2
XI18963 bl<27> cbl<13> in1<121> in2<121> sl<27> vdd vss wl<121> / cell_PIM2
XI18962 bl<27> cbl<13> in1<122> in2<122> sl<27> vdd vss wl<122> / cell_PIM2
XI17656 bl<5> cbl<2> in1<38> in2<38> sl<5> vdd vss wl<38> / cell_PIM2
XI17655 bl<5> cbl<2> in1<37> in2<37> sl<5> vdd vss wl<37> / cell_PIM2
XI17654 bl<5> cbl<2> in1<36> in2<36> sl<5> vdd vss wl<36> / cell_PIM2
XI18308 bl<13> cbl<6> in1<63> in2<63> sl<13> vdd vss wl<63> / cell_PIM2
XI18956 bl<25> cbl<12> in1<118> in2<118> sl<25> vdd vss wl<118> / cell_PIM2
XI18955 bl<25> cbl<12> in1<119> in2<119> sl<25> vdd vss wl<119> / cell_PIM2
XI18954 bl<25> cbl<12> in1<120> in2<120> sl<25> vdd vss wl<120> / cell_PIM2
XI17653 bl<5> cbl<2> in1<35> in2<35> sl<5> vdd vss wl<35> / cell_PIM2
XI17652 bl<5> cbl<2> in1<34> in2<34> sl<5> vdd vss wl<34> / cell_PIM2
XI18302 bl<11> cbl<5> in1<63> in2<63> sl<11> vdd vss wl<63> / cell_PIM2
XI18301 bl<11> cbl<5> in1<64> in2<64> sl<11> vdd vss wl<64> / cell_PIM2
XI18300 bl<11> cbl<5> in1<65> in2<65> sl<11> vdd vss wl<65> / cell_PIM2
XI18299 bl<11> cbl<5> in1<66> in2<66> sl<11> vdd vss wl<66> / cell_PIM2
XI18953 bl<25> cbl<12> in1<121> in2<121> sl<25> vdd vss wl<121> / cell_PIM2
XI18952 bl<25> cbl<12> in1<122> in2<122> sl<25> vdd vss wl<122> / cell_PIM2
XI18946 bl<23> cbl<11> in1<118> in2<118> sl<23> vdd vss wl<118> / cell_PIM2
XI18945 bl<23> cbl<11> in1<119> in2<119> sl<23> vdd vss wl<119> / cell_PIM2
XI18944 bl<23> cbl<11> in1<120> in2<120> sl<23> vdd vss wl<120> / cell_PIM2
XI18298 bl<11> cbl<5> in1<67> in2<67> sl<11> vdd vss wl<67> / cell_PIM2
XI17646 bl<7> cbl<3> in1<39> in2<39> sl<7> vdd vss wl<39> / cell_PIM2
XI17645 bl<7> cbl<3> in1<40> in2<40> sl<7> vdd vss wl<40> / cell_PIM2
XI17644 bl<7> cbl<3> in1<41> in2<41> sl<7> vdd vss wl<41> / cell_PIM2
XI17643 bl<7> cbl<3> in1<42> in2<42> sl<7> vdd vss wl<42> / cell_PIM2
XI17642 bl<7> cbl<3> in1<43> in2<43> sl<7> vdd vss wl<43> / cell_PIM2
XI18292 bl<9> cbl<4> in1<67> in2<67> sl<9> vdd vss wl<67> / cell_PIM2
XI18291 bl<9> cbl<4> in1<66> in2<66> sl<9> vdd vss wl<66> / cell_PIM2
XI18290 bl<9> cbl<4> in1<65> in2<65> sl<9> vdd vss wl<65> / cell_PIM2
XI18289 bl<9> cbl<4> in1<64> in2<64> sl<9> vdd vss wl<64> / cell_PIM2
XI18943 bl<23> cbl<11> in1<121> in2<121> sl<23> vdd vss wl<121> / cell_PIM2
XI18942 bl<23> cbl<11> in1<122> in2<122> sl<23> vdd vss wl<122> / cell_PIM2
XI17636 bl<5> cbl<2> in1<43> in2<43> sl<5> vdd vss wl<43> / cell_PIM2
XI17635 bl<5> cbl<2> in1<42> in2<42> sl<5> vdd vss wl<42> / cell_PIM2
XI17634 bl<5> cbl<2> in1<41> in2<41> sl<5> vdd vss wl<41> / cell_PIM2
XI18288 bl<9> cbl<4> in1<63> in2<63> sl<9> vdd vss wl<63> / cell_PIM2
XI18936 bl<21> cbl<10> in1<119> in2<119> sl<21> vdd vss wl<119> / cell_PIM2
XI18935 bl<21> cbl<10> in1<118> in2<118> sl<21> vdd vss wl<118> / cell_PIM2
XI18934 bl<21> cbl<10> in1<122> in2<122> sl<21> vdd vss wl<122> / cell_PIM2
XI17633 bl<5> cbl<2> in1<40> in2<40> sl<5> vdd vss wl<40> / cell_PIM2
XI17632 bl<5> cbl<2> in1<39> in2<39> sl<5> vdd vss wl<39> / cell_PIM2
XI18282 bl<15> cbl<7> in1<68> in2<68> sl<15> vdd vss wl<68> / cell_PIM2
XI18281 bl<15> cbl<7> in1<69> in2<69> sl<15> vdd vss wl<69> / cell_PIM2
XI18280 bl<15> cbl<7> in1<70> in2<70> sl<15> vdd vss wl<70> / cell_PIM2
XI18279 bl<15> cbl<7> in1<71> in2<71> sl<15> vdd vss wl<71> / cell_PIM2
XI18933 bl<21> cbl<10> in1<121> in2<121> sl<21> vdd vss wl<121> / cell_PIM2
XI18932 bl<21> cbl<10> in1<120> in2<120> sl<21> vdd vss wl<120> / cell_PIM2
XI18926 bl<19> cbl<9> in1<118> in2<118> sl<19> vdd vss wl<118> / cell_PIM2
XI18925 bl<19> cbl<9> in1<119> in2<119> sl<19> vdd vss wl<119> / cell_PIM2
XI18924 bl<19> cbl<9> in1<120> in2<120> sl<19> vdd vss wl<120> / cell_PIM2
XI18274 bl<13> cbl<6> in1<71> in2<71> sl<13> vdd vss wl<71> / cell_PIM2
XI17626 bl<7> cbl<3> in1<44> in2<44> sl<7> vdd vss wl<44> / cell_PIM2
XI17625 bl<7> cbl<3> in1<45> in2<45> sl<7> vdd vss wl<45> / cell_PIM2
XI17624 bl<7> cbl<3> in1<46> in2<46> sl<7> vdd vss wl<46> / cell_PIM2
XI17623 bl<7> cbl<3> in1<47> in2<47> sl<7> vdd vss wl<47> / cell_PIM2
XI18273 bl<13> cbl<6> in1<70> in2<70> sl<13> vdd vss wl<70> / cell_PIM2
XI18272 bl<13> cbl<6> in1<69> in2<69> sl<13> vdd vss wl<69> / cell_PIM2
XI18271 bl<13> cbl<6> in1<68> in2<68> sl<13> vdd vss wl<68> / cell_PIM2
XI18923 bl<19> cbl<9> in1<121> in2<121> sl<19> vdd vss wl<121> / cell_PIM2
XI18922 bl<19> cbl<9> in1<122> in2<122> sl<19> vdd vss wl<122> / cell_PIM2
XI17618 bl<5> cbl<2> in1<47> in2<47> sl<5> vdd vss wl<47> / cell_PIM2
XI17617 bl<5> cbl<2> in1<46> in2<46> sl<5> vdd vss wl<46> / cell_PIM2
XI17616 bl<5> cbl<2> in1<45> in2<45> sl<5> vdd vss wl<45> / cell_PIM2
XI17615 bl<5> cbl<2> in1<44> in2<44> sl<5> vdd vss wl<44> / cell_PIM2
XI18266 bl<11> cbl<5> in1<68> in2<68> sl<11> vdd vss wl<68> / cell_PIM2
XI18265 bl<11> cbl<5> in1<69> in2<69> sl<11> vdd vss wl<69> / cell_PIM2
XI18264 bl<11> cbl<5> in1<70> in2<70> sl<11> vdd vss wl<70> / cell_PIM2
XI18916 bl<17> cbl<8> in1<119> in2<119> sl<17> vdd vss wl<119> / cell_PIM2
XI18915 bl<17> cbl<8> in1<118> in2<118> sl<17> vdd vss wl<118> / cell_PIM2
XI18914 bl<17> cbl<8> in1<122> in2<122> sl<17> vdd vss wl<122> / cell_PIM2
XI17610 bl<7> cbl<3> in1<48> in2<48> sl<7> vdd vss wl<48> / cell_PIM2
XI17609 bl<7> cbl<3> in1<49> in2<49> sl<7> vdd vss wl<49> / cell_PIM2
XI18263 bl<11> cbl<5> in1<71> in2<71> sl<11> vdd vss wl<71> / cell_PIM2
XI18913 bl<17> cbl<8> in1<121> in2<121> sl<17> vdd vss wl<121> / cell_PIM2
XI18912 bl<17> cbl<8> in1<120> in2<120> sl<17> vdd vss wl<120> / cell_PIM2
XI18906 bl<31> cbl<15> in1<127> in2<127> sl<31> vdd vss wl<127> / cell_PIM2
XI18905 bl<31> cbl<15> in1<126> in2<126> sl<31> vdd vss wl<126> / cell_PIM2
XI18904 bl<31> cbl<15> in1<125> in2<125> sl<31> vdd vss wl<125> / cell_PIM2
XI18258 bl<9> cbl<4> in1<71> in2<71> sl<9> vdd vss wl<71> / cell_PIM2
XI18257 bl<9> cbl<4> in1<70> in2<70> sl<9> vdd vss wl<70> / cell_PIM2
XI18256 bl<9> cbl<4> in1<69> in2<69> sl<9> vdd vss wl<69> / cell_PIM2
XI18255 bl<9> cbl<4> in1<68> in2<68> sl<9> vdd vss wl<68> / cell_PIM2
XI17608 bl<7> cbl<3> in1<50> in2<50> sl<7> vdd vss wl<50> / cell_PIM2
XI17607 bl<7> cbl<3> in1<51> in2<51> sl<7> vdd vss wl<51> / cell_PIM2
XI17606 bl<7> cbl<3> in1<52> in2<52> sl<7> vdd vss wl<52> / cell_PIM2
XI17600 bl<5> cbl<2> in1<52> in2<52> sl<5> vdd vss wl<52> / cell_PIM2
XI17599 bl<5> cbl<2> in1<51> in2<51> sl<5> vdd vss wl<51> / cell_PIM2
XI18250 bl<15> cbl<7> in1<72> in2<72> sl<15> vdd vss wl<72> / cell_PIM2
XI18249 bl<15> cbl<7> in1<73> in2<73> sl<15> vdd vss wl<73> / cell_PIM2
XI18903 bl<31> cbl<15> in1<123> in2<123> sl<31> vdd vss wl<123> / cell_PIM2
XI18902 bl<31> cbl<15> in1<124> in2<124> sl<31> vdd vss wl<124> / cell_PIM2
XI17598 bl<5> cbl<2> in1<50> in2<50> sl<5> vdd vss wl<50> / cell_PIM2
XI17597 bl<5> cbl<2> in1<49> in2<49> sl<5> vdd vss wl<49> / cell_PIM2
XI17596 bl<5> cbl<2> in1<48> in2<48> sl<5> vdd vss wl<48> / cell_PIM2
XI18248 bl<15> cbl<7> in1<74> in2<74> sl<15> vdd vss wl<74> / cell_PIM2
XI18247 bl<15> cbl<7> in1<75> in2<75> sl<15> vdd vss wl<75> / cell_PIM2
XI18246 bl<15> cbl<7> in1<76> in2<76> sl<15> vdd vss wl<76> / cell_PIM2
XI18896 bl<29> cbl<14> in1<127> in2<127> sl<29> vdd vss wl<127> / cell_PIM2
XI18895 bl<29> cbl<14> in1<126> in2<126> sl<29> vdd vss wl<126> / cell_PIM2
XI18894 bl<29> cbl<14> in1<125> in2<125> sl<29> vdd vss wl<125> / cell_PIM2
XI17590 bl<7> cbl<3> in1<53> in2<53> sl<7> vdd vss wl<53> / cell_PIM2
XI17589 bl<7> cbl<3> in1<54> in2<54> sl<7> vdd vss wl<54> / cell_PIM2
XI18240 bl<13> cbl<6> in1<76> in2<76> sl<13> vdd vss wl<76> / cell_PIM2
XI18239 bl<13> cbl<6> in1<75> in2<75> sl<13> vdd vss wl<75> / cell_PIM2
XI18893 bl<29> cbl<14> in1<124> in2<124> sl<29> vdd vss wl<124> / cell_PIM2
XI18892 bl<29> cbl<14> in1<123> in2<123> sl<29> vdd vss wl<123> / cell_PIM2
XI18886 bl<27> cbl<13> in1<127> in2<127> sl<27> vdd vss wl<127> / cell_PIM2
XI18885 bl<27> cbl<13> in1<126> in2<126> sl<27> vdd vss wl<126> / cell_PIM2
XI18884 bl<27> cbl<13> in1<125> in2<125> sl<27> vdd vss wl<125> / cell_PIM2
XI18238 bl<13> cbl<6> in1<74> in2<74> sl<13> vdd vss wl<74> / cell_PIM2
XI18237 bl<13> cbl<6> in1<73> in2<73> sl<13> vdd vss wl<73> / cell_PIM2
XI18236 bl<13> cbl<6> in1<72> in2<72> sl<13> vdd vss wl<72> / cell_PIM2
XI17588 bl<7> cbl<3> in1<55> in2<55> sl<7> vdd vss wl<55> / cell_PIM2
XI17587 bl<7> cbl<3> in1<56> in2<56> sl<7> vdd vss wl<56> / cell_PIM2
XI17586 bl<7> cbl<3> in1<57> in2<57> sl<7> vdd vss wl<57> / cell_PIM2
XI17580 bl<5> cbl<2> in1<57> in2<57> sl<5> vdd vss wl<57> / cell_PIM2
XI17579 bl<5> cbl<2> in1<56> in2<56> sl<5> vdd vss wl<56> / cell_PIM2
XI18230 bl<11> cbl<5> in1<72> in2<72> sl<11> vdd vss wl<72> / cell_PIM2
XI18229 bl<11> cbl<5> in1<73> in2<73> sl<11> vdd vss wl<73> / cell_PIM2
XI18883 bl<27> cbl<13> in1<123> in2<123> sl<27> vdd vss wl<123> / cell_PIM2
XI18882 bl<27> cbl<13> in1<124> in2<124> sl<27> vdd vss wl<124> / cell_PIM2
XI17578 bl<5> cbl<2> in1<55> in2<55> sl<5> vdd vss wl<55> / cell_PIM2
XI17577 bl<5> cbl<2> in1<54> in2<54> sl<5> vdd vss wl<54> / cell_PIM2
XI17576 bl<5> cbl<2> in1<53> in2<53> sl<5> vdd vss wl<53> / cell_PIM2
XI18228 bl<11> cbl<5> in1<74> in2<74> sl<11> vdd vss wl<74> / cell_PIM2
XI18227 bl<11> cbl<5> in1<75> in2<75> sl<11> vdd vss wl<75> / cell_PIM2
XI18226 bl<11> cbl<5> in1<76> in2<76> sl<11> vdd vss wl<76> / cell_PIM2
XI18876 bl<25> cbl<12> in1<127> in2<127> sl<25> vdd vss wl<127> / cell_PIM2
XI18875 bl<25> cbl<12> in1<126> in2<126> sl<25> vdd vss wl<126> / cell_PIM2
XI18874 bl<25> cbl<12> in1<125> in2<125> sl<25> vdd vss wl<125> / cell_PIM2
XI17570 bl<7> cbl<3> in1<58> in2<58> sl<7> vdd vss wl<58> / cell_PIM2
XI17569 bl<7> cbl<3> in1<59> in2<59> sl<7> vdd vss wl<59> / cell_PIM2
XI18220 bl<9> cbl<4> in1<76> in2<76> sl<9> vdd vss wl<76> / cell_PIM2
XI18219 bl<9> cbl<4> in1<75> in2<75> sl<9> vdd vss wl<75> / cell_PIM2
XI18873 bl<25> cbl<12> in1<123> in2<123> sl<25> vdd vss wl<123> / cell_PIM2
XI18872 bl<25> cbl<12> in1<124> in2<124> sl<25> vdd vss wl<124> / cell_PIM2
XI18866 bl<23> cbl<11> in1<127> in2<127> sl<23> vdd vss wl<127> / cell_PIM2
XI18865 bl<23> cbl<11> in1<126> in2<126> sl<23> vdd vss wl<126> / cell_PIM2
XI18864 bl<23> cbl<11> in1<125> in2<125> sl<23> vdd vss wl<125> / cell_PIM2
XI18218 bl<9> cbl<4> in1<74> in2<74> sl<9> vdd vss wl<74> / cell_PIM2
XI18217 bl<9> cbl<4> in1<73> in2<73> sl<9> vdd vss wl<73> / cell_PIM2
XI18216 bl<9> cbl<4> in1<72> in2<72> sl<9> vdd vss wl<72> / cell_PIM2
XI17568 bl<7> cbl<3> in1<60> in2<60> sl<7> vdd vss wl<60> / cell_PIM2
XI17567 bl<7> cbl<3> in1<61> in2<61> sl<7> vdd vss wl<61> / cell_PIM2
XI17566 bl<7> cbl<3> in1<62> in2<62> sl<7> vdd vss wl<62> / cell_PIM2
XI17560 bl<5> cbl<2> in1<62> in2<62> sl<5> vdd vss wl<62> / cell_PIM2
XI17559 bl<5> cbl<2> in1<61> in2<61> sl<5> vdd vss wl<61> / cell_PIM2
XI18210 bl<15> cbl<7> in1<77> in2<77> sl<15> vdd vss wl<77> / cell_PIM2
XI18209 bl<15> cbl<7> in1<78> in2<78> sl<15> vdd vss wl<78> / cell_PIM2
XI18863 bl<23> cbl<11> in1<123> in2<123> sl<23> vdd vss wl<123> / cell_PIM2
XI18862 bl<23> cbl<11> in1<124> in2<124> sl<23> vdd vss wl<124> / cell_PIM2
XI17558 bl<5> cbl<2> in1<60> in2<60> sl<5> vdd vss wl<60> / cell_PIM2
XI17557 bl<5> cbl<2> in1<59> in2<59> sl<5> vdd vss wl<59> / cell_PIM2
XI17556 bl<5> cbl<2> in1<58> in2<58> sl<5> vdd vss wl<58> / cell_PIM2
XI18208 bl<15> cbl<7> in1<79> in2<79> sl<15> vdd vss wl<79> / cell_PIM2
XI18207 bl<15> cbl<7> in1<80> in2<80> sl<15> vdd vss wl<80> / cell_PIM2
XI18206 bl<15> cbl<7> in1<81> in2<81> sl<15> vdd vss wl<81> / cell_PIM2
XI18856 bl<21> cbl<10> in1<127> in2<127> sl<21> vdd vss wl<127> / cell_PIM2
XI18855 bl<21> cbl<10> in1<126> in2<126> sl<21> vdd vss wl<126> / cell_PIM2
XI18854 bl<21> cbl<10> in1<125> in2<125> sl<21> vdd vss wl<125> / cell_PIM2
XI17550 bl<7> cbl<3> in1<63> in2<63> sl<7> vdd vss wl<63> / cell_PIM2
XI17549 bl<7> cbl<3> in1<64> in2<64> sl<7> vdd vss wl<64> / cell_PIM2
XI18200 bl<13> cbl<6> in1<81> in2<81> sl<13> vdd vss wl<81> / cell_PIM2
XI18199 bl<13> cbl<6> in1<80> in2<80> sl<13> vdd vss wl<80> / cell_PIM2
XI18853 bl<21> cbl<10> in1<124> in2<124> sl<21> vdd vss wl<124> / cell_PIM2
XI18852 bl<21> cbl<10> in1<123> in2<123> sl<21> vdd vss wl<123> / cell_PIM2
XI18846 bl<19> cbl<9> in1<127> in2<127> sl<19> vdd vss wl<127> / cell_PIM2
XI18845 bl<19> cbl<9> in1<126> in2<126> sl<19> vdd vss wl<126> / cell_PIM2
XI18844 bl<19> cbl<9> in1<125> in2<125> sl<19> vdd vss wl<125> / cell_PIM2
XI18198 bl<13> cbl<6> in1<79> in2<79> sl<13> vdd vss wl<79> / cell_PIM2
XI18197 bl<13> cbl<6> in1<78> in2<78> sl<13> vdd vss wl<78> / cell_PIM2
XI18196 bl<13> cbl<6> in1<77> in2<77> sl<13> vdd vss wl<77> / cell_PIM2
XI17548 bl<7> cbl<3> in1<65> in2<65> sl<7> vdd vss wl<65> / cell_PIM2
XI17547 bl<7> cbl<3> in1<66> in2<66> sl<7> vdd vss wl<66> / cell_PIM2
XI17546 bl<7> cbl<3> in1<67> in2<67> sl<7> vdd vss wl<67> / cell_PIM2
XI17540 bl<5> cbl<2> in1<67> in2<67> sl<5> vdd vss wl<67> / cell_PIM2
XI17539 bl<5> cbl<2> in1<66> in2<66> sl<5> vdd vss wl<66> / cell_PIM2
XI18190 bl<11> cbl<5> in1<77> in2<77> sl<11> vdd vss wl<77> / cell_PIM2
XI18189 bl<11> cbl<5> in1<78> in2<78> sl<11> vdd vss wl<78> / cell_PIM2
XI18843 bl<19> cbl<9> in1<123> in2<123> sl<19> vdd vss wl<123> / cell_PIM2
XI18842 bl<19> cbl<9> in1<124> in2<124> sl<19> vdd vss wl<124> / cell_PIM2
XI17538 bl<5> cbl<2> in1<65> in2<65> sl<5> vdd vss wl<65> / cell_PIM2
XI17537 bl<5> cbl<2> in1<64> in2<64> sl<5> vdd vss wl<64> / cell_PIM2
XI17536 bl<5> cbl<2> in1<63> in2<63> sl<5> vdd vss wl<63> / cell_PIM2
XI18188 bl<11> cbl<5> in1<79> in2<79> sl<11> vdd vss wl<79> / cell_PIM2
XI18187 bl<11> cbl<5> in1<80> in2<80> sl<11> vdd vss wl<80> / cell_PIM2
XI18186 bl<11> cbl<5> in1<81> in2<81> sl<11> vdd vss wl<81> / cell_PIM2
XI18836 bl<17> cbl<8> in1<127> in2<127> sl<17> vdd vss wl<127> / cell_PIM2
XI18835 bl<17> cbl<8> in1<126> in2<126> sl<17> vdd vss wl<126> / cell_PIM2
XI18834 bl<17> cbl<8> in1<125> in2<125> sl<17> vdd vss wl<125> / cell_PIM2
XI17530 bl<7> cbl<3> in1<68> in2<68> sl<7> vdd vss wl<68> / cell_PIM2
XI17529 bl<7> cbl<3> in1<69> in2<69> sl<7> vdd vss wl<69> / cell_PIM2
XI18180 bl<9> cbl<4> in1<81> in2<81> sl<9> vdd vss wl<81> / cell_PIM2
XI18179 bl<9> cbl<4> in1<80> in2<80> sl<9> vdd vss wl<80> / cell_PIM2
XI18833 bl<17> cbl<8> in1<124> in2<124> sl<17> vdd vss wl<124> / cell_PIM2
XI18832 bl<17> cbl<8> in1<123> in2<123> sl<17> vdd vss wl<123> / cell_PIM2
XI18826 bl<15> cbl<7> in1<0> in2<0> sl<15> vdd vss wl<0> / cell_PIM2
XI18824 bl<13> cbl<6> in1<0> in2<0> sl<13> vdd vss wl<0> / cell_PIM2
XI18178 bl<9> cbl<4> in1<79> in2<79> sl<9> vdd vss wl<79> / cell_PIM2
XI18177 bl<9> cbl<4> in1<78> in2<78> sl<9> vdd vss wl<78> / cell_PIM2
XI18176 bl<9> cbl<4> in1<77> in2<77> sl<9> vdd vss wl<77> / cell_PIM2
XI17528 bl<7> cbl<3> in1<70> in2<70> sl<7> vdd vss wl<70> / cell_PIM2
XI17527 bl<7> cbl<3> in1<71> in2<71> sl<7> vdd vss wl<71> / cell_PIM2
XI17522 bl<5> cbl<2> in1<71> in2<71> sl<5> vdd vss wl<71> / cell_PIM2
XI17521 bl<5> cbl<2> in1<70> in2<70> sl<5> vdd vss wl<70> / cell_PIM2
XI17520 bl<5> cbl<2> in1<69> in2<69> sl<5> vdd vss wl<69> / cell_PIM2
XI17519 bl<5> cbl<2> in1<68> in2<68> sl<5> vdd vss wl<68> / cell_PIM2
XI18170 bl<15> cbl<7> in1<82> in2<82> sl<15> vdd vss wl<82> / cell_PIM2
XI18169 bl<15> cbl<7> in1<83> in2<83> sl<15> vdd vss wl<83> / cell_PIM2
XI18822 bl<11> cbl<5> in1<0> in2<0> sl<11> vdd vss wl<0> / cell_PIM2
XI18820 bl<9> cbl<4> in1<0> in2<0> sl<9> vdd vss wl<0> / cell_PIM2
XI17514 bl<7> cbl<3> in1<72> in2<72> sl<7> vdd vss wl<72> / cell_PIM2
XI18168 bl<15> cbl<7> in1<84> in2<84> sl<15> vdd vss wl<84> / cell_PIM2
XI18167 bl<15> cbl<7> in1<85> in2<85> sl<15> vdd vss wl<85> / cell_PIM2
XI18166 bl<15> cbl<7> in1<86> in2<86> sl<15> vdd vss wl<86> / cell_PIM2
XI18818 bl<15> cbl<7> in1<1> in2<1> sl<15> vdd vss wl<1> / cell_PIM2
XI18817 bl<15> cbl<7> in1<4> in2<4> sl<15> vdd vss wl<4> / cell_PIM2
XI18816 bl<15> cbl<7> in1<3> in2<3> sl<15> vdd vss wl<3> / cell_PIM2
XI18815 bl<15> cbl<7> in1<2> in2<2> sl<15> vdd vss wl<2> / cell_PIM2
XI17513 bl<7> cbl<3> in1<73> in2<73> sl<7> vdd vss wl<73> / cell_PIM2
XI17512 bl<7> cbl<3> in1<74> in2<74> sl<7> vdd vss wl<74> / cell_PIM2
XI17511 bl<7> cbl<3> in1<75> in2<75> sl<7> vdd vss wl<75> / cell_PIM2
XI17510 bl<7> cbl<3> in1<76> in2<76> sl<7> vdd vss wl<76> / cell_PIM2
XI18160 bl<13> cbl<6> in1<86> in2<86> sl<13> vdd vss wl<86> / cell_PIM2
XI18159 bl<13> cbl<6> in1<85> in2<85> sl<13> vdd vss wl<85> / cell_PIM2
XI18810 bl<13> cbl<6> in1<2> in2<2> sl<13> vdd vss wl<2> / cell_PIM2
XI18809 bl<13> cbl<6> in1<3> in2<3> sl<13> vdd vss wl<3> / cell_PIM2
XI18808 bl<13> cbl<6> in1<4> in2<4> sl<13> vdd vss wl<4> / cell_PIM2
XI18807 bl<13> cbl<6> in1<1> in2<1> sl<13> vdd vss wl<1> / cell_PIM2
XI18158 bl<13> cbl<6> in1<84> in2<84> sl<13> vdd vss wl<84> / cell_PIM2
XI18157 bl<13> cbl<6> in1<83> in2<83> sl<13> vdd vss wl<83> / cell_PIM2
XI18156 bl<13> cbl<6> in1<82> in2<82> sl<13> vdd vss wl<82> / cell_PIM2
XI17504 bl<5> cbl<2> in1<76> in2<76> sl<5> vdd vss wl<76> / cell_PIM2
XI17503 bl<5> cbl<2> in1<75> in2<75> sl<5> vdd vss wl<75> / cell_PIM2
XI17502 bl<5> cbl<2> in1<74> in2<74> sl<5> vdd vss wl<74> / cell_PIM2
XI17501 bl<5> cbl<2> in1<73> in2<73> sl<5> vdd vss wl<73> / cell_PIM2
XI17500 bl<5> cbl<2> in1<72> in2<72> sl<5> vdd vss wl<72> / cell_PIM2
XI18150 bl<11> cbl<5> in1<82> in2<82> sl<11> vdd vss wl<82> / cell_PIM2
XI18149 bl<11> cbl<5> in1<83> in2<83> sl<11> vdd vss wl<83> / cell_PIM2
XI18802 bl<11> cbl<5> in1<1> in2<1> sl<11> vdd vss wl<1> / cell_PIM2
XI18801 bl<11> cbl<5> in1<4> in2<4> sl<11> vdd vss wl<4> / cell_PIM2
XI18800 bl<11> cbl<5> in1<3> in2<3> sl<11> vdd vss wl<3> / cell_PIM2
XI18799 bl<11> cbl<5> in1<2> in2<2> sl<11> vdd vss wl<2> / cell_PIM2
XI17494 bl<7> cbl<3> in1<77> in2<77> sl<7> vdd vss wl<77> / cell_PIM2
XI18148 bl<11> cbl<5> in1<84> in2<84> sl<11> vdd vss wl<84> / cell_PIM2
XI18147 bl<11> cbl<5> in1<85> in2<85> sl<11> vdd vss wl<85> / cell_PIM2
XI18146 bl<11> cbl<5> in1<86> in2<86> sl<11> vdd vss wl<86> / cell_PIM2
XI18794 bl<9> cbl<4> in1<2> in2<2> sl<9> vdd vss wl<2> / cell_PIM2
XI16971 bl<1> cbl<0> in1<64> in2<64> sl<1> vdd vss wl<64> / cell_PIM2
XI16970 bl<1> cbl<0> in1<63> in2<63> sl<1> vdd vss wl<63> / cell_PIM2
XI16968 bl<1> cbl<0> in1<61> in2<61> sl<1> vdd vss wl<61> / cell_PIM2
XI16967 bl<1> cbl<0> in1<60> in2<60> sl<1> vdd vss wl<60> / cell_PIM2
XI16965 bl<1> cbl<0> in1<58> in2<58> sl<1> vdd vss wl<58> / cell_PIM2
XI16964 bl<1> cbl<0> in1<57> in2<57> sl<1> vdd vss wl<57> / cell_PIM2
XI16962 bl<1> cbl<0> in1<55> in2<55> sl<1> vdd vss wl<55> / cell_PIM2
XI16961 bl<1> cbl<0> in1<54> in2<54> sl<1> vdd vss wl<54> / cell_PIM2
XI16959 bl<1> cbl<0> in1<52> in2<52> sl<1> vdd vss wl<52> / cell_PIM2
XI16958 bl<1> cbl<0> in1<51> in2<51> sl<1> vdd vss wl<51> / cell_PIM2
XI16956 bl<1> cbl<0> in1<49> in2<49> sl<1> vdd vss wl<49> / cell_PIM2
XI16955 bl<1> cbl<0> in1<48> in2<48> sl<1> vdd vss wl<48> / cell_PIM2
XI16953 bl<1> cbl<0> in1<46> in2<46> sl<1> vdd vss wl<46> / cell_PIM2
XI16952 bl<1> cbl<0> in1<45> in2<45> sl<1> vdd vss wl<45> / cell_PIM2
XI16950 bl<1> cbl<0> in1<43> in2<43> sl<1> vdd vss wl<43> / cell_PIM2
XI16949 bl<1> cbl<0> in1<42> in2<42> sl<1> vdd vss wl<42> / cell_PIM2
XI16947 bl<1> cbl<0> in1<40> in2<40> sl<1> vdd vss wl<40> / cell_PIM2
XI16946 bl<1> cbl<0> in1<39> in2<39> sl<1> vdd vss wl<39> / cell_PIM2
XI16944 bl<1> cbl<0> in1<37> in2<37> sl<1> vdd vss wl<37> / cell_PIM2
XI16943 bl<1> cbl<0> in1<36> in2<36> sl<1> vdd vss wl<36> / cell_PIM2
XI16941 bl<1> cbl<0> in1<34> in2<34> sl<1> vdd vss wl<34> / cell_PIM2
XI16940 bl<1> cbl<0> in1<33> in2<33> sl<1> vdd vss wl<33> / cell_PIM2
XI16938 bl<1> cbl<0> in1<31> in2<31> sl<1> vdd vss wl<31> / cell_PIM2
XI16937 bl<1> cbl<0> in1<30> in2<30> sl<1> vdd vss wl<30> / cell_PIM2
XI16935 bl<1> cbl<0> in1<28> in2<28> sl<1> vdd vss wl<28> / cell_PIM2
XI16934 bl<1> cbl<0> in1<27> in2<27> sl<1> vdd vss wl<27> / cell_PIM2
XI16932 bl<1> cbl<0> in1<25> in2<25> sl<1> vdd vss wl<25> / cell_PIM2
XI16931 bl<1> cbl<0> in1<24> in2<24> sl<1> vdd vss wl<24> / cell_PIM2
XI16929 bl<1> cbl<0> in1<22> in2<22> sl<1> vdd vss wl<22> / cell_PIM2
XI16928 bl<1> cbl<0> in1<21> in2<21> sl<1> vdd vss wl<21> / cell_PIM2
XI16926 bl<1> cbl<0> in1<19> in2<19> sl<1> vdd vss wl<19> / cell_PIM2
XI16925 bl<1> cbl<0> in1<18> in2<18> sl<1> vdd vss wl<18> / cell_PIM2
XI16923 bl<1> cbl<0> in1<16> in2<16> sl<1> vdd vss wl<16> / cell_PIM2
XI16922 bl<1> cbl<0> in1<15> in2<15> sl<1> vdd vss wl<15> / cell_PIM2
XI16920 bl<1> cbl<0> in1<13> in2<13> sl<1> vdd vss wl<13> / cell_PIM2
XI16919 bl<1> cbl<0> in1<12> in2<12> sl<1> vdd vss wl<12> / cell_PIM2
XI16917 bl<1> cbl<0> in1<10> in2<10> sl<1> vdd vss wl<10> / cell_PIM2
XI16916 bl<1> cbl<0> in1<9> in2<9> sl<1> vdd vss wl<9> / cell_PIM2
XI16914 bl<1> cbl<0> in1<7> in2<7> sl<1> vdd vss wl<7> / cell_PIM2
XI16913 bl<1> cbl<0> in1<6> in2<6> sl<1> vdd vss wl<6> / cell_PIM2
XI16911 bl<1> cbl<0> in1<4> in2<4> sl<1> vdd vss wl<4> / cell_PIM2
XI16910 bl<1> cbl<0> in1<3> in2<3> sl<1> vdd vss wl<3> / cell_PIM2
XI16907 bl<1> cbl<0> in1<0> in2<0> sl<1> vdd vss wl<0> / cell_PIM2
XI24383 bl<61> cbl<30> in1<20> in2<20> sl<61> vdd vss wl<20> / cell_PIM2
XI25032 bl<61> cbl<30> vdd vdd sl<61> vdd vss vss / cell_PIM2
XI25030 bl<59> cbl<29> vdd vdd sl<59> vdd vss vss / cell_PIM2
XI25028 bl<57> cbl<28> vdd vdd sl<57> vdd vss vss / cell_PIM2
XI25026 bl<55> cbl<27> vdd vdd sl<55> vdd vss vss / cell_PIM2
XI25024 bl<53> cbl<26> vdd vdd sl<53> vdd vss vss / cell_PIM2
XI24378 bl<59> cbl<29> in1<18> in2<18> sl<59> vdd vss wl<18> / cell_PIM2
XI25022 bl<51> cbl<25> vdd vdd sl<51> vdd vss vss / cell_PIM2
XI25020 bl<49> cbl<24> vdd vdd sl<49> vdd vss vss / cell_PIM2
XI24368 bl<57> cbl<28> in1<20> in2<20> sl<57> vdd vss wl<20> / cell_PIM2
XI25016 bl<45> cbl<22> vdd vdd sl<45> vdd vss vss / cell_PIM2
XI25014 bl<43> cbl<21> vdd vdd sl<43> vdd vss vss / cell_PIM2
XI25018 bl<47> cbl<23> vdd vdd sl<47> vdd vss vss / cell_PIM2
XI25012 bl<41> cbl<20> vdd vdd sl<41> vdd vss vss / cell_PIM2
XI25010 bl<39> cbl<19> vdd vdd sl<39> vdd vss vss / cell_PIM2
XI25008 bl<37> cbl<18> vdd vdd sl<37> vdd vss vss / cell_PIM2
XI25006 bl<35> cbl<17> vdd vdd sl<35> vdd vss vss / cell_PIM2
XI25004 bl<33> cbl<16> vdd vdd sl<33> vdd vss vss / cell_PIM2
XI24353 bl<53> cbl<26> in1<18> in2<18> sl<53> vdd vss wl<18> / cell_PIM2
XI25002 bl<31> cbl<15> vdd vdd sl<31> vdd vss vss / cell_PIM2
XI25000 bl<29> cbl<14> vdd vdd sl<29> vdd vss vss / cell_PIM2
XI24996 bl<25> cbl<12> vdd vdd sl<25> vdd vss vss / cell_PIM2
XI24994 bl<23> cbl<11> vdd vdd sl<23> vdd vss vss / cell_PIM2
XI24998 bl<27> cbl<13> vdd vdd sl<27> vdd vss vss / cell_PIM2
XI24343 bl<51> cbl<25> in1<21> in2<21> sl<51> vdd vss wl<21> / cell_PIM2
XI24992 bl<21> cbl<10> vdd vdd sl<21> vdd vss vss / cell_PIM2
XI24990 bl<19> cbl<9> vdd vdd sl<19> vdd vss vss / cell_PIM2
XI24988 bl<17> cbl<8> vdd vdd sl<17> vdd vss vss / cell_PIM2
XI24986 bl<15> cbl<7> vdd vdd sl<15> vdd vss vss / cell_PIM2
XI24984 bl<13> cbl<6> vdd vdd sl<13> vdd vss vss / cell_PIM2
XI24338 bl<49> cbl<24> in1<19> in2<19> sl<49> vdd vss wl<19> / cell_PIM2
XI24982 bl<11> cbl<5> vdd vdd sl<11> vdd vss vss / cell_PIM2
XI24980 bl<9> cbl<4> vdd vdd sl<9> vdd vss vss / cell_PIM2
XI24328 bl<47> cbl<23> in1<20> in2<20> sl<47> vdd vss wl<20> / cell_PIM2
XI24976 bl<5> cbl<2> vdd vdd sl<5> vdd vss vss / cell_PIM2
XI24974 bl<3> cbl<1> vdd vdd sl<3> vdd vss vss / cell_PIM2
XI24978 bl<7> cbl<3> vdd vdd sl<7> vdd vss vss / cell_PIM2
XI24972 bl<1> cbl<0> vdd vdd sl<1> vdd vss vss / cell_PIM2
XI24970 bl<63> cbl<31> in1<0> in2<0> sl<63> vdd vss wl<0> / cell_PIM2
XI24969 bl<63> cbl<31> in1<1> in2<1> sl<63> vdd vss wl<1> / cell_PIM2
XI24968 bl<63> cbl<31> in1<2> in2<2> sl<63> vdd vss wl<2> / cell_PIM2
XI24964 bl<61> cbl<30> in1<0> in2<0> sl<61> vdd vss wl<0> / cell_PIM2
XI24313 bl<43> cbl<21> in1<19> in2<19> sl<43> vdd vss wl<19> / cell_PIM2
XI24962 bl<61> cbl<30> in1<1> in2<1> sl<61> vdd vss wl<1> / cell_PIM2
XI24963 bl<61> cbl<30> in1<2> in2<2> sl<61> vdd vss wl<2> / cell_PIM2
XI24957 bl<59> cbl<29> in1<1> in2<1> sl<59> vdd vss wl<1> / cell_PIM2
XI24956 bl<59> cbl<29> in1<2> in2<2> sl<59> vdd vss wl<2> / cell_PIM2
XI24958 bl<59> cbl<29> in1<0> in2<0> sl<59> vdd vss wl<0> / cell_PIM2
XI24303 bl<41> cbl<20> in1<21> in2<21> sl<41> vdd vss wl<21> / cell_PIM2
XI24952 bl<57> cbl<28> in1<0> in2<0> sl<57> vdd vss wl<0> / cell_PIM2
XI24951 bl<57> cbl<28> in1<1> in2<1> sl<57> vdd vss wl<1> / cell_PIM2
XI24950 bl<57> cbl<28> in1<2> in2<2> sl<57> vdd vss wl<2> / cell_PIM2
XI24946 bl<55> cbl<27> in1<0> in2<0> sl<55> vdd vss wl<0> / cell_PIM2
XI24945 bl<55> cbl<27> in1<1> in2<1> sl<55> vdd vss wl<1> / cell_PIM2
XI24944 bl<55> cbl<27> in1<2> in2<2> sl<55> vdd vss wl<2> / cell_PIM2
XI24298 bl<39> cbl<19> in1<18> in2<18> sl<39> vdd vss wl<18> / cell_PIM2
XI24940 bl<53> cbl<26> in1<0> in2<0> sl<53> vdd vss wl<0> / cell_PIM2
XI24939 bl<53> cbl<26> in1<2> in2<2> sl<53> vdd vss wl<2> / cell_PIM2
XI24288 bl<37> cbl<18> in1<21> in2<21> sl<37> vdd vss wl<21> / cell_PIM2
XI24934 bl<51> cbl<25> in1<0> in2<0> sl<51> vdd vss wl<0> / cell_PIM2
XI24938 bl<53> cbl<26> in1<1> in2<1> sl<53> vdd vss wl<1> / cell_PIM2
XI24932 bl<51> cbl<25> in1<2> in2<2> sl<51> vdd vss wl<2> / cell_PIM2
XI24933 bl<51> cbl<25> in1<1> in2<1> sl<51> vdd vss wl<1> / cell_PIM2
XI24928 bl<49> cbl<24> in1<0> in2<0> sl<49> vdd vss wl<0> / cell_PIM2
XI24927 bl<49> cbl<24> in1<2> in2<2> sl<49> vdd vss wl<2> / cell_PIM2
XI24926 bl<49> cbl<24> in1<1> in2<1> sl<49> vdd vss wl<1> / cell_PIM2
XI24273 bl<33> cbl<16> in1<18> in2<18> sl<33> vdd vss wl<18> / cell_PIM2
XI24922 bl<47> cbl<23> in1<0> in2<0> sl<47> vdd vss wl<0> / cell_PIM2
XI24921 bl<47> cbl<23> in1<1> in2<1> sl<47> vdd vss wl<1> / cell_PIM2
XI24920 bl<47> cbl<23> in1<2> in2<2> sl<47> vdd vss wl<2> / cell_PIM2
XI24916 bl<45> cbl<22> in1<0> in2<0> sl<45> vdd vss wl<0> / cell_PIM2
XI24915 bl<45> cbl<22> in1<2> in2<2> sl<45> vdd vss wl<2> / cell_PIM2
XI24914 bl<45> cbl<22> in1<1> in2<1> sl<45> vdd vss wl<1> / cell_PIM2
XI24263 bl<63> cbl<31> in1<25> in2<25> sl<63> vdd vss wl<25> / cell_PIM2
XI24910 bl<43> cbl<21> in1<0> in2<0> sl<43> vdd vss wl<0> / cell_PIM2
XI24909 bl<43> cbl<21> in1<1> in2<1> sl<43> vdd vss wl<1> / cell_PIM2
XI24908 bl<43> cbl<21> in1<2> in2<2> sl<43> vdd vss wl<2> / cell_PIM2
XI24904 bl<41> cbl<20> in1<0> in2<0> sl<41> vdd vss wl<0> / cell_PIM2
XI24253 bl<61> cbl<30> in1<26> in2<26> sl<61> vdd vss wl<26> / cell_PIM2
XI24902 bl<41> cbl<20> in1<2> in2<2> sl<41> vdd vss wl<2> / cell_PIM2
XI24903 bl<41> cbl<20> in1<1> in2<1> sl<41> vdd vss wl<1> / cell_PIM2
XI24897 bl<39> cbl<19> in1<1> in2<1> sl<39> vdd vss wl<1> / cell_PIM2
XI24896 bl<39> cbl<19> in1<2> in2<2> sl<39> vdd vss wl<2> / cell_PIM2
XI24898 bl<39> cbl<19> in1<0> in2<0> sl<39> vdd vss wl<0> / cell_PIM2
XI24243 bl<59> cbl<29> in1<25> in2<25> sl<59> vdd vss wl<25> / cell_PIM2
XI24892 bl<37> cbl<18> in1<0> in2<0> sl<37> vdd vss wl<0> / cell_PIM2
XI24891 bl<37> cbl<18> in1<2> in2<2> sl<37> vdd vss wl<2> / cell_PIM2
XI24890 bl<37> cbl<18> in1<1> in2<1> sl<37> vdd vss wl<1> / cell_PIM2
XI24886 bl<35> cbl<17> in1<0> in2<0> sl<35> vdd vss wl<0> / cell_PIM2
XI24885 bl<35> cbl<17> in1<1> in2<1> sl<35> vdd vss wl<1> / cell_PIM2
XI24884 bl<35> cbl<17> in1<2> in2<2> sl<35> vdd vss wl<2> / cell_PIM2
XI24233 bl<57> cbl<28> in1<25> in2<25> sl<57> vdd vss wl<25> / cell_PIM2
XI24880 bl<33> cbl<16> in1<0> in2<0> sl<33> vdd vss wl<0> / cell_PIM2
XI24879 bl<33> cbl<16> in1<2> in2<2> sl<33> vdd vss wl<2> / cell_PIM2
XI24874 bl<63> cbl<31> in1<4> in2<4> sl<63> vdd vss wl<4> / cell_PIM2
XI24878 bl<33> cbl<16> in1<1> in2<1> sl<33> vdd vss wl<1> / cell_PIM2
XI23148 bl<57> cbl<28> in1<56> in2<56> sl<57> vdd vss wl<56> / cell_PIM2
XI23147 bl<57> cbl<28> in1<57> in2<57> sl<57> vdd vss wl<57> / cell_PIM2
XI23146 bl<57> cbl<28> in1<58> in2<58> sl<57> vdd vss wl<58> / cell_PIM2
XI23145 bl<57> cbl<28> in1<59> in2<59> sl<57> vdd vss wl<59> / cell_PIM2
XI23730 bl<49> cbl<24> in1<38> in2<38> sl<49> vdd vss wl<38> / cell_PIM2
XI23729 bl<49> cbl<24> in1<37> in2<37> sl<49> vdd vss wl<37> / cell_PIM2
XI24377 bl<59> cbl<29> in1<19> in2<19> sl<59> vdd vss wl<19> / cell_PIM2
XI24376 bl<59> cbl<29> in1<20> in2<20> sl<59> vdd vss wl<20> / cell_PIM2
XI24375 bl<59> cbl<29> in1<21> in2<21> sl<59> vdd vss wl<21> / cell_PIM2
XI23728 bl<49> cbl<24> in1<40> in2<40> sl<49> vdd vss wl<40> / cell_PIM2
XI23727 bl<49> cbl<24> in1<39> in2<39> sl<49> vdd vss wl<39> / cell_PIM2
XI23144 bl<57> cbl<28> in1<60> in2<60> sl<57> vdd vss wl<60> / cell_PIM2
XI22558 bl<61> cbl<30> in1<79> in2<79> sl<61> vdd vss wl<79> / cell_PIM2
XI23138 bl<55> cbl<27> in1<56> in2<56> sl<55> vdd vss wl<56> / cell_PIM2
XI23137 bl<55> cbl<27> in1<57> in2<57> sl<55> vdd vss wl<57> / cell_PIM2
XI23722 bl<47> cbl<23> in1<37> in2<37> sl<47> vdd vss wl<37> / cell_PIM2
XI23721 bl<47> cbl<23> in1<38> in2<38> sl<47> vdd vss wl<38> / cell_PIM2
XI23720 bl<47> cbl<23> in1<39> in2<39> sl<47> vdd vss wl<39> / cell_PIM2
XI23719 bl<47> cbl<23> in1<40> in2<40> sl<47> vdd vss wl<40> / cell_PIM2
XI24370 bl<57> cbl<28> in1<18> in2<18> sl<57> vdd vss wl<18> / cell_PIM2
XI24369 bl<57> cbl<28> in1<19> in2<19> sl<57> vdd vss wl<19> / cell_PIM2
XI22548 bl<59> cbl<29> in1<77> in2<77> sl<59> vdd vss wl<77> / cell_PIM2
XI23136 bl<55> cbl<27> in1<58> in2<58> sl<55> vdd vss wl<58> / cell_PIM2
XI23135 bl<55> cbl<27> in1<59> in2<59> sl<55> vdd vss wl<59> / cell_PIM2
XI23134 bl<55> cbl<27> in1<60> in2<60> sl<55> vdd vss wl<60> / cell_PIM2
XI23714 bl<45> cbl<22> in1<38> in2<38> sl<45> vdd vss wl<38> / cell_PIM2
XI24367 bl<57> cbl<28> in1<21> in2<21> sl<57> vdd vss wl<21> / cell_PIM2
XI23713 bl<45> cbl<22> in1<37> in2<37> sl<45> vdd vss wl<37> / cell_PIM2
XI23712 bl<45> cbl<22> in1<40> in2<40> sl<45> vdd vss wl<40> / cell_PIM2
XI23711 bl<45> cbl<22> in1<39> in2<39> sl<45> vdd vss wl<39> / cell_PIM2
XI24362 bl<55> cbl<27> in1<18> in2<18> sl<55> vdd vss wl<18> / cell_PIM2
XI24361 bl<55> cbl<27> in1<19> in2<19> sl<55> vdd vss wl<19> / cell_PIM2
XI24360 bl<55> cbl<27> in1<20> in2<20> sl<55> vdd vss wl<20> / cell_PIM2
XI24359 bl<55> cbl<27> in1<21> in2<21> sl<55> vdd vss wl<21> / cell_PIM2
XI24354 bl<53> cbl<26> in1<19> in2<19> sl<53> vdd vss wl<19> / cell_PIM2
XI23706 bl<43> cbl<21> in1<37> in2<37> sl<43> vdd vss wl<37> / cell_PIM2
XI23705 bl<43> cbl<21> in1<38> in2<38> sl<43> vdd vss wl<38> / cell_PIM2
XI23704 bl<43> cbl<21> in1<39> in2<39> sl<43> vdd vss wl<39> / cell_PIM2
XI23128 bl<53> cbl<26> in1<57> in2<57> sl<53> vdd vss wl<57> / cell_PIM2
XI23127 bl<53> cbl<26> in1<56> in2<56> sl<53> vdd vss wl<56> / cell_PIM2
XI23126 bl<53> cbl<26> in1<60> in2<60> sl<53> vdd vss wl<60> / cell_PIM2
XI23125 bl<53> cbl<26> in1<59> in2<59> sl<53> vdd vss wl<59> / cell_PIM2
XI22538 bl<57> cbl<28> in1<77> in2<77> sl<57> vdd vss wl<77> / cell_PIM2
XI23124 bl<53> cbl<26> in1<58> in2<58> sl<53> vdd vss wl<58> / cell_PIM2
XI23703 bl<43> cbl<21> in1<40> in2<40> sl<43> vdd vss wl<40> / cell_PIM2
XI24352 bl<53> cbl<26> in1<21> in2<21> sl<53> vdd vss wl<21> / cell_PIM2
XI24351 bl<53> cbl<26> in1<20> in2<20> sl<53> vdd vss wl<20> / cell_PIM2
XI22528 bl<55> cbl<27> in1<77> in2<77> sl<55> vdd vss wl<77> / cell_PIM2
XI23118 bl<51> cbl<25> in1<56> in2<56> sl<51> vdd vss wl<56> / cell_PIM2
XI23117 bl<51> cbl<25> in1<57> in2<57> sl<51> vdd vss wl<57> / cell_PIM2
XI23698 bl<41> cbl<20> in1<37> in2<37> sl<41> vdd vss wl<37> / cell_PIM2
XI23697 bl<41> cbl<20> in1<38> in2<38> sl<41> vdd vss wl<38> / cell_PIM2
XI23696 bl<41> cbl<20> in1<39> in2<39> sl<41> vdd vss wl<39> / cell_PIM2
XI23695 bl<41> cbl<20> in1<40> in2<40> sl<41> vdd vss wl<40> / cell_PIM2
XI24346 bl<51> cbl<25> in1<18> in2<18> sl<51> vdd vss wl<18> / cell_PIM2
XI24345 bl<51> cbl<25> in1<19> in2<19> sl<51> vdd vss wl<19> / cell_PIM2
XI24344 bl<51> cbl<25> in1<20> in2<20> sl<51> vdd vss wl<20> / cell_PIM2
XI23116 bl<51> cbl<25> in1<58> in2<58> sl<51> vdd vss wl<58> / cell_PIM2
XI23115 bl<51> cbl<25> in1<59> in2<59> sl<51> vdd vss wl<59> / cell_PIM2
XI23114 bl<51> cbl<25> in1<60> in2<60> sl<51> vdd vss wl<60> / cell_PIM2
XI23690 bl<39> cbl<19> in1<37> in2<37> sl<39> vdd vss wl<37> / cell_PIM2
XI23689 bl<39> cbl<19> in1<38> in2<38> sl<39> vdd vss wl<38> / cell_PIM2
XI24337 bl<49> cbl<24> in1<18> in2<18> sl<49> vdd vss wl<18> / cell_PIM2
XI24336 bl<49> cbl<24> in1<21> in2<21> sl<49> vdd vss wl<21> / cell_PIM2
XI24335 bl<49> cbl<24> in1<20> in2<20> sl<49> vdd vss wl<20> / cell_PIM2
XI23688 bl<39> cbl<19> in1<39> in2<39> sl<39> vdd vss wl<39> / cell_PIM2
XI23687 bl<39> cbl<19> in1<40> in2<40> sl<39> vdd vss wl<40> / cell_PIM2
XI22518 bl<53> cbl<26> in1<79> in2<79> sl<53> vdd vss wl<79> / cell_PIM2
XI23108 bl<49> cbl<24> in1<57> in2<57> sl<49> vdd vss wl<57> / cell_PIM2
XI23107 bl<49> cbl<24> in1<56> in2<56> sl<49> vdd vss wl<56> / cell_PIM2
XI23106 bl<49> cbl<24> in1<60> in2<60> sl<49> vdd vss wl<60> / cell_PIM2
XI23105 bl<49> cbl<24> in1<59> in2<59> sl<49> vdd vss wl<59> / cell_PIM2
XI23682 bl<37> cbl<18> in1<38> in2<38> sl<37> vdd vss wl<38> / cell_PIM2
XI23681 bl<37> cbl<18> in1<37> in2<37> sl<37> vdd vss wl<37> / cell_PIM2
XI23680 bl<37> cbl<18> in1<40> in2<40> sl<37> vdd vss wl<40> / cell_PIM2
XI23679 bl<37> cbl<18> in1<39> in2<39> sl<37> vdd vss wl<39> / cell_PIM2
XI24330 bl<47> cbl<23> in1<18> in2<18> sl<47> vdd vss wl<18> / cell_PIM2
XI24329 bl<47> cbl<23> in1<19> in2<19> sl<47> vdd vss wl<19> / cell_PIM2
XI22508 bl<51> cbl<25> in1<77> in2<77> sl<51> vdd vss wl<77> / cell_PIM2
XI23104 bl<49> cbl<24> in1<58> in2<58> sl<49> vdd vss wl<58> / cell_PIM2
XI23674 bl<35> cbl<17> in1<37> in2<37> sl<35> vdd vss wl<37> / cell_PIM2
XI24327 bl<47> cbl<23> in1<21> in2<21> sl<47> vdd vss wl<21> / cell_PIM2
XI23098 bl<47> cbl<23> in1<56> in2<56> sl<47> vdd vss wl<56> / cell_PIM2
XI23097 bl<47> cbl<23> in1<57> in2<57> sl<47> vdd vss wl<57> / cell_PIM2
XI23673 bl<35> cbl<17> in1<38> in2<38> sl<35> vdd vss wl<38> / cell_PIM2
XI23672 bl<35> cbl<17> in1<39> in2<39> sl<35> vdd vss wl<39> / cell_PIM2
XI23671 bl<35> cbl<17> in1<40> in2<40> sl<35> vdd vss wl<40> / cell_PIM2
XI24322 bl<45> cbl<22> in1<19> in2<19> sl<45> vdd vss wl<19> / cell_PIM2
XI24321 bl<45> cbl<22> in1<18> in2<18> sl<45> vdd vss wl<18> / cell_PIM2
XI24320 bl<45> cbl<22> in1<21> in2<21> sl<45> vdd vss wl<21> / cell_PIM2
XI24319 bl<45> cbl<22> in1<20> in2<20> sl<45> vdd vss wl<20> / cell_PIM2
XI24314 bl<43> cbl<21> in1<18> in2<18> sl<43> vdd vss wl<18> / cell_PIM2
XI23666 bl<33> cbl<16> in1<38> in2<38> sl<33> vdd vss wl<38> / cell_PIM2
XI23665 bl<33> cbl<16> in1<37> in2<37> sl<33> vdd vss wl<37> / cell_PIM2
XI23664 bl<33> cbl<16> in1<40> in2<40> sl<33> vdd vss wl<40> / cell_PIM2
XI23096 bl<47> cbl<23> in1<58> in2<58> sl<47> vdd vss wl<58> / cell_PIM2
XI23095 bl<47> cbl<23> in1<59> in2<59> sl<47> vdd vss wl<59> / cell_PIM2
XI23094 bl<47> cbl<23> in1<60> in2<60> sl<47> vdd vss wl<60> / cell_PIM2
XI22498 bl<49> cbl<24> in1<79> in2<79> sl<49> vdd vss wl<79> / cell_PIM2
XI23663 bl<33> cbl<16> in1<39> in2<39> sl<33> vdd vss wl<39> / cell_PIM2
XI24312 bl<43> cbl<21> in1<20> in2<20> sl<43> vdd vss wl<20> / cell_PIM2
XI24311 bl<43> cbl<21> in1<21> in2<21> sl<43> vdd vss wl<21> / cell_PIM2
XI22488 bl<47> cbl<23> in1<77> in2<77> sl<47> vdd vss wl<77> / cell_PIM2
XI23088 bl<45> cbl<22> in1<57> in2<57> sl<45> vdd vss wl<57> / cell_PIM2
XI23087 bl<45> cbl<22> in1<56> in2<56> sl<45> vdd vss wl<56> / cell_PIM2
XI23086 bl<45> cbl<22> in1<60> in2<60> sl<45> vdd vss wl<60> / cell_PIM2
XI23085 bl<45> cbl<22> in1<59> in2<59> sl<45> vdd vss wl<59> / cell_PIM2
XI23658 bl<63> cbl<31> in1<41> in2<41> sl<63> vdd vss wl<41> / cell_PIM2
XI23657 bl<63> cbl<31> in1<42> in2<42> sl<63> vdd vss wl<42> / cell_PIM2
XI23656 bl<63> cbl<31> in1<43> in2<43> sl<63> vdd vss wl<43> / cell_PIM2
XI23655 bl<63> cbl<31> in1<44> in2<44> sl<63> vdd vss wl<44> / cell_PIM2
XI23654 bl<63> cbl<31> in1<45> in2<45> sl<63> vdd vss wl<45> / cell_PIM2
XI24306 bl<41> cbl<20> in1<18> in2<18> sl<41> vdd vss wl<18> / cell_PIM2
XI24305 bl<41> cbl<20> in1<19> in2<19> sl<41> vdd vss wl<19> / cell_PIM2
XI24304 bl<41> cbl<20> in1<20> in2<20> sl<41> vdd vss wl<20> / cell_PIM2
XI23084 bl<45> cbl<22> in1<58> in2<58> sl<45> vdd vss wl<58> / cell_PIM2
XI24297 bl<39> cbl<19> in1<19> in2<19> sl<39> vdd vss wl<19> / cell_PIM2
XI24296 bl<39> cbl<19> in1<20> in2<20> sl<39> vdd vss wl<20> / cell_PIM2
XI24295 bl<39> cbl<19> in1<21> in2<21> sl<39> vdd vss wl<21> / cell_PIM2
XI23648 bl<61> cbl<30> in1<43> in2<43> sl<61> vdd vss wl<43> / cell_PIM2
XI23647 bl<61> cbl<30> in1<42> in2<42> sl<61> vdd vss wl<42> / cell_PIM2
XI23646 bl<61> cbl<30> in1<41> in2<41> sl<61> vdd vss wl<41> / cell_PIM2
XI23645 bl<61> cbl<30> in1<45> in2<45> sl<61> vdd vss wl<45> / cell_PIM2
XI23644 bl<61> cbl<30> in1<44> in2<44> sl<61> vdd vss wl<44> / cell_PIM2
XI23078 bl<43> cbl<21> in1<56> in2<56> sl<43> vdd vss wl<56> / cell_PIM2
XI23077 bl<43> cbl<21> in1<57> in2<57> sl<43> vdd vss wl<57> / cell_PIM2
XI22478 bl<45> cbl<22> in1<79> in2<79> sl<45> vdd vss wl<79> / cell_PIM2
XI23076 bl<43> cbl<21> in1<58> in2<58> sl<43> vdd vss wl<58> / cell_PIM2
XI23075 bl<43> cbl<21> in1<59> in2<59> sl<43> vdd vss wl<59> / cell_PIM2
XI23074 bl<43> cbl<21> in1<60> in2<60> sl<43> vdd vss wl<60> / cell_PIM2
XI24290 bl<37> cbl<18> in1<19> in2<19> sl<37> vdd vss wl<19> / cell_PIM2
XI24289 bl<37> cbl<18> in1<18> in2<18> sl<37> vdd vss wl<18> / cell_PIM2
XI22468 bl<43> cbl<21> in1<77> in2<77> sl<43> vdd vss wl<77> / cell_PIM2
XI23638 bl<59> cbl<29> in1<41> in2<41> sl<59> vdd vss wl<41> / cell_PIM2
XI23637 bl<59> cbl<29> in1<42> in2<42> sl<59> vdd vss wl<42> / cell_PIM2
XI23636 bl<59> cbl<29> in1<43> in2<43> sl<59> vdd vss wl<43> / cell_PIM2
XI23635 bl<59> cbl<29> in1<44> in2<44> sl<59> vdd vss wl<44> / cell_PIM2
XI23634 bl<59> cbl<29> in1<45> in2<45> sl<59> vdd vss wl<45> / cell_PIM2
XI24287 bl<37> cbl<18> in1<20> in2<20> sl<37> vdd vss wl<20> / cell_PIM2
XI23068 bl<41> cbl<20> in1<56> in2<56> sl<41> vdd vss wl<56> / cell_PIM2
XI23067 bl<41> cbl<20> in1<57> in2<57> sl<41> vdd vss wl<57> / cell_PIM2
XI23066 bl<41> cbl<20> in1<58> in2<58> sl<41> vdd vss wl<58> / cell_PIM2
XI23065 bl<41> cbl<20> in1<59> in2<59> sl<41> vdd vss wl<59> / cell_PIM2
XI24282 bl<35> cbl<17> in1<18> in2<18> sl<35> vdd vss wl<18> / cell_PIM2
XI24281 bl<35> cbl<17> in1<19> in2<19> sl<35> vdd vss wl<19> / cell_PIM2
XI24280 bl<35> cbl<17> in1<20> in2<20> sl<35> vdd vss wl<20> / cell_PIM2
XI24279 bl<35> cbl<17> in1<21> in2<21> sl<35> vdd vss wl<21> / cell_PIM2
XI24274 bl<33> cbl<16> in1<19> in2<19> sl<33> vdd vss wl<19> / cell_PIM2
XI23628 bl<57> cbl<28> in1<41> in2<41> sl<57> vdd vss wl<41> / cell_PIM2
XI23627 bl<57> cbl<28> in1<42> in2<42> sl<57> vdd vss wl<42> / cell_PIM2
XI23626 bl<57> cbl<28> in1<43> in2<43> sl<57> vdd vss wl<43> / cell_PIM2
XI23625 bl<57> cbl<28> in1<44> in2<44> sl<57> vdd vss wl<44> / cell_PIM2
XI23624 bl<57> cbl<28> in1<45> in2<45> sl<57> vdd vss wl<45> / cell_PIM2
XI23064 bl<41> cbl<20> in1<60> in2<60> sl<41> vdd vss wl<60> / cell_PIM2
XI22458 bl<41> cbl<20> in1<77> in2<77> sl<41> vdd vss wl<77> / cell_PIM2
XI23058 bl<39> cbl<19> in1<56> in2<56> sl<39> vdd vss wl<56> / cell_PIM2
XI23057 bl<39> cbl<19> in1<57> in2<57> sl<39> vdd vss wl<57> / cell_PIM2
XI24272 bl<33> cbl<16> in1<21> in2<21> sl<33> vdd vss wl<21> / cell_PIM2
XI24271 bl<33> cbl<16> in1<20> in2<20> sl<33> vdd vss wl<20> / cell_PIM2
XI22448 bl<39> cbl<19> in1<77> in2<77> sl<39> vdd vss wl<77> / cell_PIM2
XI23056 bl<39> cbl<19> in1<58> in2<58> sl<39> vdd vss wl<58> / cell_PIM2
XI23055 bl<39> cbl<19> in1<59> in2<59> sl<39> vdd vss wl<59> / cell_PIM2
XI23054 bl<39> cbl<19> in1<60> in2<60> sl<39> vdd vss wl<60> / cell_PIM2
XI23618 bl<55> cbl<27> in1<41> in2<41> sl<55> vdd vss wl<41> / cell_PIM2
XI23617 bl<55> cbl<27> in1<42> in2<42> sl<55> vdd vss wl<42> / cell_PIM2
XI23616 bl<55> cbl<27> in1<43> in2<43> sl<55> vdd vss wl<43> / cell_PIM2
XI23615 bl<55> cbl<27> in1<44> in2<44> sl<55> vdd vss wl<44> / cell_PIM2
XI23614 bl<55> cbl<27> in1<45> in2<45> sl<55> vdd vss wl<45> / cell_PIM2
XI24266 bl<63> cbl<31> in1<22> in2<22> sl<63> vdd vss wl<22> / cell_PIM2
XI24265 bl<63> cbl<31> in1<23> in2<23> sl<63> vdd vss wl<23> / cell_PIM2
XI24264 bl<63> cbl<31> in1<24> in2<24> sl<63> vdd vss wl<24> / cell_PIM2
XI24262 bl<63> cbl<31> in1<26> in2<26> sl<63> vdd vss wl<26> / cell_PIM2
XI24256 bl<61> cbl<30> in1<24> in2<24> sl<61> vdd vss wl<24> / cell_PIM2
XI24255 bl<61> cbl<30> in1<23> in2<23> sl<61> vdd vss wl<23> / cell_PIM2
XI24254 bl<61> cbl<30> in1<22> in2<22> sl<61> vdd vss wl<22> / cell_PIM2
XI23608 bl<53> cbl<26> in1<43> in2<43> sl<53> vdd vss wl<43> / cell_PIM2
XI23607 bl<53> cbl<26> in1<42> in2<42> sl<53> vdd vss wl<42> / cell_PIM2
XI23606 bl<53> cbl<26> in1<41> in2<41> sl<53> vdd vss wl<41> / cell_PIM2
XI23605 bl<53> cbl<26> in1<45> in2<45> sl<53> vdd vss wl<45> / cell_PIM2
XI23604 bl<53> cbl<26> in1<44> in2<44> sl<53> vdd vss wl<44> / cell_PIM2
XI23048 bl<37> cbl<18> in1<57> in2<57> sl<37> vdd vss wl<57> / cell_PIM2
XI23047 bl<37> cbl<18> in1<56> in2<56> sl<37> vdd vss wl<56> / cell_PIM2
XI23046 bl<37> cbl<18> in1<60> in2<60> sl<37> vdd vss wl<60> / cell_PIM2
XI23045 bl<37> cbl<18> in1<59> in2<59> sl<37> vdd vss wl<59> / cell_PIM2
XI22438 bl<37> cbl<18> in1<79> in2<79> sl<37> vdd vss wl<79> / cell_PIM2
XI23044 bl<37> cbl<18> in1<58> in2<58> sl<37> vdd vss wl<58> / cell_PIM2
XI24252 bl<61> cbl<30> in1<25> in2<25> sl<61> vdd vss wl<25> / cell_PIM2
XI22428 bl<35> cbl<17> in1<77> in2<77> sl<35> vdd vss wl<77> / cell_PIM2
XI23038 bl<35> cbl<17> in1<56> in2<56> sl<35> vdd vss wl<56> / cell_PIM2
XI23037 bl<35> cbl<17> in1<57> in2<57> sl<35> vdd vss wl<57> / cell_PIM2
XI23598 bl<51> cbl<25> in1<41> in2<41> sl<51> vdd vss wl<41> / cell_PIM2
XI23597 bl<51> cbl<25> in1<42> in2<42> sl<51> vdd vss wl<42> / cell_PIM2
XI23596 bl<51> cbl<25> in1<43> in2<43> sl<51> vdd vss wl<43> / cell_PIM2
XI23595 bl<51> cbl<25> in1<44> in2<44> sl<51> vdd vss wl<44> / cell_PIM2
XI23594 bl<51> cbl<25> in1<45> in2<45> sl<51> vdd vss wl<45> / cell_PIM2
XI24246 bl<59> cbl<29> in1<22> in2<22> sl<59> vdd vss wl<22> / cell_PIM2
XI24245 bl<59> cbl<29> in1<23> in2<23> sl<59> vdd vss wl<23> / cell_PIM2
XI24244 bl<59> cbl<29> in1<24> in2<24> sl<59> vdd vss wl<24> / cell_PIM2
XI23036 bl<35> cbl<17> in1<58> in2<58> sl<35> vdd vss wl<58> / cell_PIM2
XI23035 bl<35> cbl<17> in1<59> in2<59> sl<35> vdd vss wl<59> / cell_PIM2
XI23034 bl<35> cbl<17> in1<60> in2<60> sl<35> vdd vss wl<60> / cell_PIM2
XI24242 bl<59> cbl<29> in1<26> in2<26> sl<59> vdd vss wl<26> / cell_PIM2
XI24236 bl<57> cbl<28> in1<22> in2<22> sl<57> vdd vss wl<22> / cell_PIM2
XI24235 bl<57> cbl<28> in1<23> in2<23> sl<57> vdd vss wl<23> / cell_PIM2
XI24234 bl<57> cbl<28> in1<24> in2<24> sl<57> vdd vss wl<24> / cell_PIM2
XI23588 bl<49> cbl<24> in1<43> in2<43> sl<49> vdd vss wl<43> / cell_PIM2
XI23587 bl<49> cbl<24> in1<42> in2<42> sl<49> vdd vss wl<42> / cell_PIM2
XI23586 bl<49> cbl<24> in1<41> in2<41> sl<49> vdd vss wl<41> / cell_PIM2
XI23585 bl<49> cbl<24> in1<45> in2<45> sl<49> vdd vss wl<45> / cell_PIM2
XI23584 bl<49> cbl<24> in1<44> in2<44> sl<49> vdd vss wl<44> / cell_PIM2
XI22418 bl<33> cbl<16> in1<79> in2<79> sl<33> vdd vss wl<79> / cell_PIM2
XI23028 bl<33> cbl<16> in1<57> in2<57> sl<33> vdd vss wl<57> / cell_PIM2
XI23027 bl<33> cbl<16> in1<56> in2<56> sl<33> vdd vss wl<56> / cell_PIM2
XI23026 bl<33> cbl<16> in1<60> in2<60> sl<33> vdd vss wl<60> / cell_PIM2
XI23025 bl<33> cbl<16> in1<59> in2<59> sl<33> vdd vss wl<59> / cell_PIM2
XI24232 bl<57> cbl<28> in1<26> in2<26> sl<57> vdd vss wl<26> / cell_PIM2
XI22408 bl<63> cbl<31> in1<82> in2<82> sl<63> vdd vss wl<82> / cell_PIM2
XI23024 bl<33> cbl<16> in1<58> in2<58> sl<33> vdd vss wl<58> / cell_PIM2
XI23578 bl<47> cbl<23> in1<41> in2<41> sl<47> vdd vss wl<41> / cell_PIM2
XI23577 bl<47> cbl<23> in1<42> in2<42> sl<47> vdd vss wl<42> / cell_PIM2
XI23576 bl<47> cbl<23> in1<43> in2<43> sl<47> vdd vss wl<43> / cell_PIM2
XI23575 bl<47> cbl<23> in1<44> in2<44> sl<47> vdd vss wl<44> / cell_PIM2
XI23574 bl<47> cbl<23> in1<45> in2<45> sl<47> vdd vss wl<45> / cell_PIM2
XI24226 bl<55> cbl<27> in1<22> in2<22> sl<55> vdd vss wl<22> / cell_PIM2
XI24225 bl<55> cbl<27> in1<23> in2<23> sl<55> vdd vss wl<23> / cell_PIM2
XI24224 bl<55> cbl<27> in1<24> in2<24> sl<55> vdd vss wl<24> / cell_PIM2
XI21263 bl<45> cbl<22> in1<114> in2<114> sl<45> vdd vss wl<114> / cell_PIM2
XI21262 bl<45> cbl<22> in1<113> in2<113> sl<45> vdd vss wl<113> / cell_PIM2
XI21261 bl<45> cbl<22> in1<117> in2<117> sl<45> vdd vss wl<117> / cell_PIM2
XI21260 bl<45> cbl<22> in1<116> in2<116> sl<45> vdd vss wl<116> / cell_PIM2
XI21912 bl<53> cbl<26> in1<95> in2<95> sl<53> vdd vss wl<95> / cell_PIM2
XI21911 bl<53> cbl<26> in1<94> in2<94> sl<53> vdd vss wl<94> / cell_PIM2
XI21910 bl<53> cbl<26> in1<98> in2<98> sl<53> vdd vss wl<98> / cell_PIM2
XI21909 bl<53> cbl<26> in1<97> in2<97> sl<53> vdd vss wl<97> / cell_PIM2
XI22560 bl<61> cbl<30> in1<76> in2<76> sl<61> vdd vss wl<76> / cell_PIM2
XI22559 bl<61> cbl<30> in1<75> in2<75> sl<61> vdd vss wl<75> / cell_PIM2
XI22557 bl<61> cbl<30> in1<78> in2<78> sl<61> vdd vss wl<78> / cell_PIM2
XI22556 bl<61> cbl<30> in1<77> in2<77> sl<61> vdd vss wl<77> / cell_PIM2
XI21908 bl<53> cbl<26> in1<96> in2<96> sl<53> vdd vss wl<96> / cell_PIM2
XI21254 bl<43> cbl<21> in1<113> in2<113> sl<43> vdd vss wl<113> / cell_PIM2
XI21253 bl<43> cbl<21> in1<114> in2<114> sl<43> vdd vss wl<114> / cell_PIM2
XI21252 bl<43> cbl<21> in1<115> in2<115> sl<43> vdd vss wl<115> / cell_PIM2
XI21251 bl<43> cbl<21> in1<116> in2<116> sl<43> vdd vss wl<116> / cell_PIM2
XI21250 bl<43> cbl<21> in1<117> in2<117> sl<43> vdd vss wl<117> / cell_PIM2
XI21902 bl<51> cbl<25> in1<94> in2<94> sl<51> vdd vss wl<94> / cell_PIM2
XI21901 bl<51> cbl<25> in1<95> in2<95> sl<51> vdd vss wl<95> / cell_PIM2
XI21900 bl<51> cbl<25> in1<96> in2<96> sl<51> vdd vss wl<96> / cell_PIM2
XI21899 bl<51> cbl<25> in1<97> in2<97> sl<51> vdd vss wl<97> / cell_PIM2
XI22550 bl<59> cbl<29> in1<75> in2<75> sl<59> vdd vss wl<75> / cell_PIM2
XI22549 bl<59> cbl<29> in1<76> in2<76> sl<59> vdd vss wl<76> / cell_PIM2
XI21244 bl<41> cbl<20> in1<113> in2<113> sl<41> vdd vss wl<113> / cell_PIM2
XI21898 bl<51> cbl<25> in1<98> in2<98> sl<51> vdd vss wl<98> / cell_PIM2
XI22547 bl<59> cbl<29> in1<78> in2<78> sl<59> vdd vss wl<78> / cell_PIM2
XI22546 bl<59> cbl<29> in1<79> in2<79> sl<59> vdd vss wl<79> / cell_PIM2
XI21243 bl<41> cbl<20> in1<114> in2<114> sl<41> vdd vss wl<114> / cell_PIM2
XI21242 bl<41> cbl<20> in1<115> in2<115> sl<41> vdd vss wl<115> / cell_PIM2
XI21241 bl<41> cbl<20> in1<116> in2<116> sl<41> vdd vss wl<116> / cell_PIM2
XI21240 bl<41> cbl<20> in1<117> in2<117> sl<41> vdd vss wl<117> / cell_PIM2
XI21892 bl<49> cbl<24> in1<95> in2<95> sl<49> vdd vss wl<95> / cell_PIM2
XI21891 bl<49> cbl<24> in1<94> in2<94> sl<49> vdd vss wl<94> / cell_PIM2
XI21890 bl<49> cbl<24> in1<98> in2<98> sl<49> vdd vss wl<98> / cell_PIM2
XI21889 bl<49> cbl<24> in1<97> in2<97> sl<49> vdd vss wl<97> / cell_PIM2
XI22540 bl<57> cbl<28> in1<75> in2<75> sl<57> vdd vss wl<75> / cell_PIM2
XI22539 bl<57> cbl<28> in1<76> in2<76> sl<57> vdd vss wl<76> / cell_PIM2
XI22537 bl<57> cbl<28> in1<78> in2<78> sl<57> vdd vss wl<78> / cell_PIM2
XI22536 bl<57> cbl<28> in1<79> in2<79> sl<57> vdd vss wl<79> / cell_PIM2
XI21888 bl<49> cbl<24> in1<96> in2<96> sl<49> vdd vss wl<96> / cell_PIM2
XI21234 bl<39> cbl<19> in1<113> in2<113> sl<39> vdd vss wl<113> / cell_PIM2
XI21233 bl<39> cbl<19> in1<114> in2<114> sl<39> vdd vss wl<114> / cell_PIM2
XI21232 bl<39> cbl<19> in1<115> in2<115> sl<39> vdd vss wl<115> / cell_PIM2
XI21231 bl<39> cbl<19> in1<116> in2<116> sl<39> vdd vss wl<116> / cell_PIM2
XI21230 bl<39> cbl<19> in1<117> in2<117> sl<39> vdd vss wl<117> / cell_PIM2
XI21882 bl<47> cbl<23> in1<94> in2<94> sl<47> vdd vss wl<94> / cell_PIM2
XI21881 bl<47> cbl<23> in1<95> in2<95> sl<47> vdd vss wl<95> / cell_PIM2
XI21880 bl<47> cbl<23> in1<96> in2<96> sl<47> vdd vss wl<96> / cell_PIM2
XI21879 bl<47> cbl<23> in1<97> in2<97> sl<47> vdd vss wl<97> / cell_PIM2
XI22530 bl<55> cbl<27> in1<75> in2<75> sl<55> vdd vss wl<75> / cell_PIM2
XI22529 bl<55> cbl<27> in1<76> in2<76> sl<55> vdd vss wl<76> / cell_PIM2
XI21224 bl<37> cbl<18> in1<115> in2<115> sl<37> vdd vss wl<115> / cell_PIM2
XI21878 bl<47> cbl<23> in1<98> in2<98> sl<47> vdd vss wl<98> / cell_PIM2
XI22527 bl<55> cbl<27> in1<78> in2<78> sl<55> vdd vss wl<78> / cell_PIM2
XI22526 bl<55> cbl<27> in1<79> in2<79> sl<55> vdd vss wl<79> / cell_PIM2
XI21223 bl<37> cbl<18> in1<114> in2<114> sl<37> vdd vss wl<114> / cell_PIM2
XI21222 bl<37> cbl<18> in1<113> in2<113> sl<37> vdd vss wl<113> / cell_PIM2
XI21221 bl<37> cbl<18> in1<117> in2<117> sl<37> vdd vss wl<117> / cell_PIM2
XI21220 bl<37> cbl<18> in1<116> in2<116> sl<37> vdd vss wl<116> / cell_PIM2
XI21872 bl<45> cbl<22> in1<95> in2<95> sl<45> vdd vss wl<95> / cell_PIM2
XI21871 bl<45> cbl<22> in1<94> in2<94> sl<45> vdd vss wl<94> / cell_PIM2
XI21870 bl<45> cbl<22> in1<98> in2<98> sl<45> vdd vss wl<98> / cell_PIM2
XI21869 bl<45> cbl<22> in1<97> in2<97> sl<45> vdd vss wl<97> / cell_PIM2
XI22520 bl<53> cbl<26> in1<76> in2<76> sl<53> vdd vss wl<76> / cell_PIM2
XI22519 bl<53> cbl<26> in1<75> in2<75> sl<53> vdd vss wl<75> / cell_PIM2
XI22517 bl<53> cbl<26> in1<78> in2<78> sl<53> vdd vss wl<78> / cell_PIM2
XI22516 bl<53> cbl<26> in1<77> in2<77> sl<53> vdd vss wl<77> / cell_PIM2
XI21868 bl<45> cbl<22> in1<96> in2<96> sl<45> vdd vss wl<96> / cell_PIM2
XI21214 bl<35> cbl<17> in1<113> in2<113> sl<35> vdd vss wl<113> / cell_PIM2
XI21213 bl<35> cbl<17> in1<114> in2<114> sl<35> vdd vss wl<114> / cell_PIM2
XI21212 bl<35> cbl<17> in1<115> in2<115> sl<35> vdd vss wl<115> / cell_PIM2
XI21211 bl<35> cbl<17> in1<116> in2<116> sl<35> vdd vss wl<116> / cell_PIM2
XI21210 bl<35> cbl<17> in1<117> in2<117> sl<35> vdd vss wl<117> / cell_PIM2
XI21862 bl<43> cbl<21> in1<94> in2<94> sl<43> vdd vss wl<94> / cell_PIM2
XI21861 bl<43> cbl<21> in1<95> in2<95> sl<43> vdd vss wl<95> / cell_PIM2
XI21860 bl<43> cbl<21> in1<96> in2<96> sl<43> vdd vss wl<96> / cell_PIM2
XI21859 bl<43> cbl<21> in1<97> in2<97> sl<43> vdd vss wl<97> / cell_PIM2
XI22510 bl<51> cbl<25> in1<75> in2<75> sl<51> vdd vss wl<75> / cell_PIM2
XI22509 bl<51> cbl<25> in1<76> in2<76> sl<51> vdd vss wl<76> / cell_PIM2
XI21204 bl<33> cbl<16> in1<115> in2<115> sl<33> vdd vss wl<115> / cell_PIM2
XI21858 bl<43> cbl<21> in1<98> in2<98> sl<43> vdd vss wl<98> / cell_PIM2
XI22507 bl<51> cbl<25> in1<78> in2<78> sl<51> vdd vss wl<78> / cell_PIM2
XI22506 bl<51> cbl<25> in1<79> in2<79> sl<51> vdd vss wl<79> / cell_PIM2
XI21203 bl<33> cbl<16> in1<114> in2<114> sl<33> vdd vss wl<114> / cell_PIM2
XI21202 bl<33> cbl<16> in1<113> in2<113> sl<33> vdd vss wl<113> / cell_PIM2
XI21201 bl<33> cbl<16> in1<117> in2<117> sl<33> vdd vss wl<117> / cell_PIM2
XI21200 bl<33> cbl<16> in1<116> in2<116> sl<33> vdd vss wl<116> / cell_PIM2
XI21852 bl<41> cbl<20> in1<94> in2<94> sl<41> vdd vss wl<94> / cell_PIM2
XI21851 bl<41> cbl<20> in1<95> in2<95> sl<41> vdd vss wl<95> / cell_PIM2
XI21850 bl<41> cbl<20> in1<96> in2<96> sl<41> vdd vss wl<96> / cell_PIM2
XI21849 bl<41> cbl<20> in1<97> in2<97> sl<41> vdd vss wl<97> / cell_PIM2
XI22500 bl<49> cbl<24> in1<76> in2<76> sl<49> vdd vss wl<76> / cell_PIM2
XI22499 bl<49> cbl<24> in1<75> in2<75> sl<49> vdd vss wl<75> / cell_PIM2
XI22497 bl<49> cbl<24> in1<78> in2<78> sl<49> vdd vss wl<78> / cell_PIM2
XI22496 bl<49> cbl<24> in1<77> in2<77> sl<49> vdd vss wl<77> / cell_PIM2
XI21848 bl<41> cbl<20> in1<98> in2<98> sl<41> vdd vss wl<98> / cell_PIM2
XI21194 bl<63> cbl<31> in1<118> in2<118> sl<63> vdd vss wl<118> / cell_PIM2
XI21193 bl<63> cbl<31> in1<119> in2<119> sl<63> vdd vss wl<119> / cell_PIM2
XI21192 bl<63> cbl<31> in1<120> in2<120> sl<63> vdd vss wl<120> / cell_PIM2
XI21191 bl<63> cbl<31> in1<121> in2<121> sl<63> vdd vss wl<121> / cell_PIM2
XI21190 bl<63> cbl<31> in1<122> in2<122> sl<63> vdd vss wl<122> / cell_PIM2
XI21842 bl<39> cbl<19> in1<94> in2<94> sl<39> vdd vss wl<94> / cell_PIM2
XI21841 bl<39> cbl<19> in1<95> in2<95> sl<39> vdd vss wl<95> / cell_PIM2
XI21840 bl<39> cbl<19> in1<96> in2<96> sl<39> vdd vss wl<96> / cell_PIM2
XI21839 bl<39> cbl<19> in1<97> in2<97> sl<39> vdd vss wl<97> / cell_PIM2
XI22490 bl<47> cbl<23> in1<75> in2<75> sl<47> vdd vss wl<75> / cell_PIM2
XI22489 bl<47> cbl<23> in1<76> in2<76> sl<47> vdd vss wl<76> / cell_PIM2
XI21184 bl<61> cbl<30> in1<119> in2<119> sl<61> vdd vss wl<119> / cell_PIM2
XI21838 bl<39> cbl<19> in1<98> in2<98> sl<39> vdd vss wl<98> / cell_PIM2
XI22487 bl<47> cbl<23> in1<78> in2<78> sl<47> vdd vss wl<78> / cell_PIM2
XI22486 bl<47> cbl<23> in1<79> in2<79> sl<47> vdd vss wl<79> / cell_PIM2
XI21183 bl<61> cbl<30> in1<118> in2<118> sl<61> vdd vss wl<118> / cell_PIM2
XI21182 bl<61> cbl<30> in1<122> in2<122> sl<61> vdd vss wl<122> / cell_PIM2
XI21181 bl<61> cbl<30> in1<121> in2<121> sl<61> vdd vss wl<121> / cell_PIM2
XI21180 bl<61> cbl<30> in1<120> in2<120> sl<61> vdd vss wl<120> / cell_PIM2
XI21832 bl<37> cbl<18> in1<95> in2<95> sl<37> vdd vss wl<95> / cell_PIM2
XI21831 bl<37> cbl<18> in1<94> in2<94> sl<37> vdd vss wl<94> / cell_PIM2
XI21830 bl<37> cbl<18> in1<98> in2<98> sl<37> vdd vss wl<98> / cell_PIM2
XI21829 bl<37> cbl<18> in1<97> in2<97> sl<37> vdd vss wl<97> / cell_PIM2
XI22480 bl<45> cbl<22> in1<76> in2<76> sl<45> vdd vss wl<76> / cell_PIM2
XI22479 bl<45> cbl<22> in1<75> in2<75> sl<45> vdd vss wl<75> / cell_PIM2
XI22477 bl<45> cbl<22> in1<78> in2<78> sl<45> vdd vss wl<78> / cell_PIM2
XI22476 bl<45> cbl<22> in1<77> in2<77> sl<45> vdd vss wl<77> / cell_PIM2
XI21828 bl<37> cbl<18> in1<96> in2<96> sl<37> vdd vss wl<96> / cell_PIM2
XI21174 bl<59> cbl<29> in1<118> in2<118> sl<59> vdd vss wl<118> / cell_PIM2
XI21173 bl<59> cbl<29> in1<119> in2<119> sl<59> vdd vss wl<119> / cell_PIM2
XI21172 bl<59> cbl<29> in1<120> in2<120> sl<59> vdd vss wl<120> / cell_PIM2
XI21171 bl<59> cbl<29> in1<121> in2<121> sl<59> vdd vss wl<121> / cell_PIM2
XI21170 bl<59> cbl<29> in1<122> in2<122> sl<59> vdd vss wl<122> / cell_PIM2
XI21822 bl<35> cbl<17> in1<94> in2<94> sl<35> vdd vss wl<94> / cell_PIM2
XI21821 bl<35> cbl<17> in1<95> in2<95> sl<35> vdd vss wl<95> / cell_PIM2
XI21820 bl<35> cbl<17> in1<96> in2<96> sl<35> vdd vss wl<96> / cell_PIM2
XI21819 bl<35> cbl<17> in1<97> in2<97> sl<35> vdd vss wl<97> / cell_PIM2
XI22470 bl<43> cbl<21> in1<75> in2<75> sl<43> vdd vss wl<75> / cell_PIM2
XI22469 bl<43> cbl<21> in1<76> in2<76> sl<43> vdd vss wl<76> / cell_PIM2
XI21164 bl<57> cbl<28> in1<118> in2<118> sl<57> vdd vss wl<118> / cell_PIM2
XI21818 bl<35> cbl<17> in1<98> in2<98> sl<35> vdd vss wl<98> / cell_PIM2
XI22467 bl<43> cbl<21> in1<78> in2<78> sl<43> vdd vss wl<78> / cell_PIM2
XI22466 bl<43> cbl<21> in1<79> in2<79> sl<43> vdd vss wl<79> / cell_PIM2
XI21163 bl<57> cbl<28> in1<119> in2<119> sl<57> vdd vss wl<119> / cell_PIM2
XI21162 bl<57> cbl<28> in1<120> in2<120> sl<57> vdd vss wl<120> / cell_PIM2
XI21161 bl<57> cbl<28> in1<121> in2<121> sl<57> vdd vss wl<121> / cell_PIM2
XI21160 bl<57> cbl<28> in1<122> in2<122> sl<57> vdd vss wl<122> / cell_PIM2
XI21812 bl<33> cbl<16> in1<95> in2<95> sl<33> vdd vss wl<95> / cell_PIM2
XI21811 bl<33> cbl<16> in1<94> in2<94> sl<33> vdd vss wl<94> / cell_PIM2
XI21810 bl<33> cbl<16> in1<98> in2<98> sl<33> vdd vss wl<98> / cell_PIM2
XI21809 bl<33> cbl<16> in1<97> in2<97> sl<33> vdd vss wl<97> / cell_PIM2
XI22460 bl<41> cbl<20> in1<75> in2<75> sl<41> vdd vss wl<75> / cell_PIM2
XI22459 bl<41> cbl<20> in1<76> in2<76> sl<41> vdd vss wl<76> / cell_PIM2
XI22457 bl<41> cbl<20> in1<78> in2<78> sl<41> vdd vss wl<78> / cell_PIM2
XI22456 bl<41> cbl<20> in1<79> in2<79> sl<41> vdd vss wl<79> / cell_PIM2
XI21808 bl<33> cbl<16> in1<96> in2<96> sl<33> vdd vss wl<96> / cell_PIM2
XI21154 bl<55> cbl<27> in1<118> in2<118> sl<55> vdd vss wl<118> / cell_PIM2
XI21153 bl<55> cbl<27> in1<119> in2<119> sl<55> vdd vss wl<119> / cell_PIM2
XI21152 bl<55> cbl<27> in1<120> in2<120> sl<55> vdd vss wl<120> / cell_PIM2
XI21151 bl<55> cbl<27> in1<121> in2<121> sl<55> vdd vss wl<121> / cell_PIM2
XI21150 bl<55> cbl<27> in1<122> in2<122> sl<55> vdd vss wl<122> / cell_PIM2
XI21802 bl<63> cbl<31> in1<99> in2<99> sl<63> vdd vss wl<99> / cell_PIM2
XI21801 bl<63> cbl<31> in1<100> in2<100> sl<63> vdd vss wl<100> / cell_PIM2
XI21800 bl<63> cbl<31> in1<101> in2<101> sl<63> vdd vss wl<101> / cell_PIM2
XI21799 bl<63> cbl<31> in1<102> in2<102> sl<63> vdd vss wl<102> / cell_PIM2
XI22450 bl<39> cbl<19> in1<75> in2<75> sl<39> vdd vss wl<75> / cell_PIM2
XI22449 bl<39> cbl<19> in1<76> in2<76> sl<39> vdd vss wl<76> / cell_PIM2
XI21144 bl<53> cbl<26> in1<119> in2<119> sl<53> vdd vss wl<119> / cell_PIM2
XI21798 bl<63> cbl<31> in1<103> in2<103> sl<63> vdd vss wl<103> / cell_PIM2
XI22447 bl<39> cbl<19> in1<78> in2<78> sl<39> vdd vss wl<78> / cell_PIM2
XI22446 bl<39> cbl<19> in1<79> in2<79> sl<39> vdd vss wl<79> / cell_PIM2
XI21143 bl<53> cbl<26> in1<118> in2<118> sl<53> vdd vss wl<118> / cell_PIM2
XI21142 bl<53> cbl<26> in1<122> in2<122> sl<53> vdd vss wl<122> / cell_PIM2
XI21141 bl<53> cbl<26> in1<121> in2<121> sl<53> vdd vss wl<121> / cell_PIM2
XI21140 bl<53> cbl<26> in1<120> in2<120> sl<53> vdd vss wl<120> / cell_PIM2
XI21792 bl<61> cbl<30> in1<100> in2<100> sl<61> vdd vss wl<100> / cell_PIM2
XI21791 bl<61> cbl<30> in1<99> in2<99> sl<61> vdd vss wl<99> / cell_PIM2
XI21790 bl<61> cbl<30> in1<103> in2<103> sl<61> vdd vss wl<103> / cell_PIM2
XI21789 bl<61> cbl<30> in1<102> in2<102> sl<61> vdd vss wl<102> / cell_PIM2
XI22440 bl<37> cbl<18> in1<76> in2<76> sl<37> vdd vss wl<76> / cell_PIM2
XI22439 bl<37> cbl<18> in1<75> in2<75> sl<37> vdd vss wl<75> / cell_PIM2
XI22437 bl<37> cbl<18> in1<78> in2<78> sl<37> vdd vss wl<78> / cell_PIM2
XI22436 bl<37> cbl<18> in1<77> in2<77> sl<37> vdd vss wl<77> / cell_PIM2
XI21788 bl<61> cbl<30> in1<101> in2<101> sl<61> vdd vss wl<101> / cell_PIM2
XI21134 bl<51> cbl<25> in1<118> in2<118> sl<51> vdd vss wl<118> / cell_PIM2
XI21133 bl<51> cbl<25> in1<119> in2<119> sl<51> vdd vss wl<119> / cell_PIM2
XI21132 bl<51> cbl<25> in1<120> in2<120> sl<51> vdd vss wl<120> / cell_PIM2
XI21131 bl<51> cbl<25> in1<121> in2<121> sl<51> vdd vss wl<121> / cell_PIM2
XI21130 bl<51> cbl<25> in1<122> in2<122> sl<51> vdd vss wl<122> / cell_PIM2
XI21782 bl<59> cbl<29> in1<99> in2<99> sl<59> vdd vss wl<99> / cell_PIM2
XI21781 bl<59> cbl<29> in1<100> in2<100> sl<59> vdd vss wl<100> / cell_PIM2
XI21780 bl<59> cbl<29> in1<101> in2<101> sl<59> vdd vss wl<101> / cell_PIM2
XI21779 bl<59> cbl<29> in1<102> in2<102> sl<59> vdd vss wl<102> / cell_PIM2
XI22430 bl<35> cbl<17> in1<75> in2<75> sl<35> vdd vss wl<75> / cell_PIM2
XI22429 bl<35> cbl<17> in1<76> in2<76> sl<35> vdd vss wl<76> / cell_PIM2
XI21124 bl<49> cbl<24> in1<119> in2<119> sl<49> vdd vss wl<119> / cell_PIM2
XI21778 bl<59> cbl<29> in1<103> in2<103> sl<59> vdd vss wl<103> / cell_PIM2
XI22427 bl<35> cbl<17> in1<78> in2<78> sl<35> vdd vss wl<78> / cell_PIM2
XI22426 bl<35> cbl<17> in1<79> in2<79> sl<35> vdd vss wl<79> / cell_PIM2
XI21123 bl<49> cbl<24> in1<118> in2<118> sl<49> vdd vss wl<118> / cell_PIM2
XI21122 bl<49> cbl<24> in1<122> in2<122> sl<49> vdd vss wl<122> / cell_PIM2
XI21121 bl<49> cbl<24> in1<121> in2<121> sl<49> vdd vss wl<121> / cell_PIM2
XI21120 bl<49> cbl<24> in1<120> in2<120> sl<49> vdd vss wl<120> / cell_PIM2
XI21772 bl<57> cbl<28> in1<99> in2<99> sl<57> vdd vss wl<99> / cell_PIM2
XI21771 bl<57> cbl<28> in1<100> in2<100> sl<57> vdd vss wl<100> / cell_PIM2
XI21770 bl<57> cbl<28> in1<101> in2<101> sl<57> vdd vss wl<101> / cell_PIM2
XI21769 bl<57> cbl<28> in1<102> in2<102> sl<57> vdd vss wl<102> / cell_PIM2
XI22420 bl<33> cbl<16> in1<76> in2<76> sl<33> vdd vss wl<76> / cell_PIM2
XI22419 bl<33> cbl<16> in1<75> in2<75> sl<33> vdd vss wl<75> / cell_PIM2
XI22417 bl<33> cbl<16> in1<78> in2<78> sl<33> vdd vss wl<78> / cell_PIM2
XI22416 bl<33> cbl<16> in1<77> in2<77> sl<33> vdd vss wl<77> / cell_PIM2
XI21768 bl<57> cbl<28> in1<103> in2<103> sl<57> vdd vss wl<103> / cell_PIM2
XI21114 bl<47> cbl<23> in1<118> in2<118> sl<47> vdd vss wl<118> / cell_PIM2
XI21113 bl<47> cbl<23> in1<119> in2<119> sl<47> vdd vss wl<119> / cell_PIM2
XI21112 bl<47> cbl<23> in1<120> in2<120> sl<47> vdd vss wl<120> / cell_PIM2
XI21111 bl<47> cbl<23> in1<121> in2<121> sl<47> vdd vss wl<121> / cell_PIM2
XI21110 bl<47> cbl<23> in1<122> in2<122> sl<47> vdd vss wl<122> / cell_PIM2
XI21762 bl<55> cbl<27> in1<99> in2<99> sl<55> vdd vss wl<99> / cell_PIM2
XI21761 bl<55> cbl<27> in1<100> in2<100> sl<55> vdd vss wl<100> / cell_PIM2
XI21760 bl<55> cbl<27> in1<101> in2<101> sl<55> vdd vss wl<101> / cell_PIM2
XI21759 bl<55> cbl<27> in1<102> in2<102> sl<55> vdd vss wl<102> / cell_PIM2
XI22410 bl<63> cbl<31> in1<80> in2<80> sl<63> vdd vss wl<80> / cell_PIM2
XI22409 bl<63> cbl<31> in1<81> in2<81> sl<63> vdd vss wl<81> / cell_PIM2
XI21104 bl<45> cbl<22> in1<119> in2<119> sl<45> vdd vss wl<119> / cell_PIM2
XI21758 bl<55> cbl<27> in1<103> in2<103> sl<55> vdd vss wl<103> / cell_PIM2
XI22407 bl<63> cbl<31> in1<83> in2<83> sl<63> vdd vss wl<83> / cell_PIM2
XI19440 bl<29> cbl<14> in1<91> in2<91> sl<29> vdd vss wl<91> / cell_PIM2
XI19439 bl<29> cbl<14> in1<90> in2<90> sl<29> vdd vss wl<90> / cell_PIM2
XI20028 bl<25> cbl<12> in1<51> in2<51> sl<25> vdd vss wl<51> / cell_PIM2
XI20027 bl<25> cbl<12> in1<52> in2<52> sl<25> vdd vss wl<52> / cell_PIM2
XI20026 bl<25> cbl<12> in1<53> in2<53> sl<25> vdd vss wl<53> / cell_PIM2
XI20025 bl<25> cbl<12> in1<54> in2<54> sl<25> vdd vss wl<54> / cell_PIM2
XI20613 bl<21> cbl<10> in1<16> in2<16> sl<21> vdd vss wl<16> / cell_PIM2
XI20612 bl<21> cbl<10> in1<15> in2<15> sl<21> vdd vss wl<15> / cell_PIM2
XI20606 bl<19> cbl<9> in1<13> in2<13> sl<19> vdd vss wl<13> / cell_PIM2
XI20605 bl<19> cbl<9> in1<14> in2<14> sl<19> vdd vss wl<14> / cell_PIM2
XI20604 bl<19> cbl<9> in1<15> in2<15> sl<19> vdd vss wl<15> / cell_PIM2
XI20024 bl<25> cbl<12> in1<55> in2<55> sl<25> vdd vss wl<55> / cell_PIM2
XI19438 bl<29> cbl<14> in1<89> in2<89> sl<29> vdd vss wl<89> / cell_PIM2
XI19437 bl<29> cbl<14> in1<93> in2<93> sl<29> vdd vss wl<93> / cell_PIM2
XI19436 bl<29> cbl<14> in1<92> in2<92> sl<29> vdd vss wl<92> / cell_PIM2
XI19430 bl<27> cbl<13> in1<89> in2<89> sl<27> vdd vss wl<89> / cell_PIM2
XI19429 bl<27> cbl<13> in1<90> in2<90> sl<27> vdd vss wl<90> / cell_PIM2
XI20018 bl<23> cbl<11> in1<51> in2<51> sl<23> vdd vss wl<51> / cell_PIM2
XI20017 bl<23> cbl<11> in1<52> in2<52> sl<23> vdd vss wl<52> / cell_PIM2
XI20603 bl<19> cbl<9> in1<16> in2<16> sl<19> vdd vss wl<16> / cell_PIM2
XI20602 bl<19> cbl<9> in1<17> in2<17> sl<19> vdd vss wl<17> / cell_PIM2
XI19427 bl<27> cbl<13> in1<92> in2<92> sl<27> vdd vss wl<92> / cell_PIM2
XI19426 bl<27> cbl<13> in1<93> in2<93> sl<27> vdd vss wl<93> / cell_PIM2
XI19428 bl<27> cbl<13> in1<91> in2<91> sl<27> vdd vss wl<91> / cell_PIM2
XI20016 bl<23> cbl<11> in1<53> in2<53> sl<23> vdd vss wl<53> / cell_PIM2
XI20015 bl<23> cbl<11> in1<54> in2<54> sl<23> vdd vss wl<54> / cell_PIM2
XI20014 bl<23> cbl<11> in1<55> in2<55> sl<23> vdd vss wl<55> / cell_PIM2
XI20596 bl<17> cbl<8> in1<14> in2<14> sl<17> vdd vss wl<14> / cell_PIM2
XI20595 bl<17> cbl<8> in1<13> in2<13> sl<17> vdd vss wl<13> / cell_PIM2
XI20594 bl<17> cbl<8> in1<17> in2<17> sl<17> vdd vss wl<17> / cell_PIM2
XI19420 bl<25> cbl<12> in1<89> in2<89> sl<25> vdd vss wl<89> / cell_PIM2
XI19419 bl<25> cbl<12> in1<90> in2<90> sl<25> vdd vss wl<90> / cell_PIM2
XI20593 bl<17> cbl<8> in1<16> in2<16> sl<17> vdd vss wl<16> / cell_PIM2
XI20592 bl<17> cbl<8> in1<15> in2<15> sl<17> vdd vss wl<15> / cell_PIM2
XI20586 bl<31> cbl<15> in1<18> in2<18> sl<31> vdd vss wl<18> / cell_PIM2
XI20585 bl<31> cbl<15> in1<19> in2<19> sl<31> vdd vss wl<19> / cell_PIM2
XI20584 bl<31> cbl<15> in1<20> in2<20> sl<31> vdd vss wl<20> / cell_PIM2
XI20008 bl<21> cbl<10> in1<52> in2<52> sl<21> vdd vss wl<52> / cell_PIM2
XI20007 bl<21> cbl<10> in1<51> in2<51> sl<21> vdd vss wl<51> / cell_PIM2
XI20006 bl<21> cbl<10> in1<55> in2<55> sl<21> vdd vss wl<55> / cell_PIM2
XI20005 bl<21> cbl<10> in1<54> in2<54> sl<21> vdd vss wl<54> / cell_PIM2
XI19418 bl<25> cbl<12> in1<91> in2<91> sl<25> vdd vss wl<91> / cell_PIM2
XI19417 bl<25> cbl<12> in1<92> in2<92> sl<25> vdd vss wl<92> / cell_PIM2
XI19416 bl<25> cbl<12> in1<93> in2<93> sl<25> vdd vss wl<93> / cell_PIM2
XI19410 bl<23> cbl<11> in1<89> in2<89> sl<23> vdd vss wl<89> / cell_PIM2
XI19409 bl<23> cbl<11> in1<90> in2<90> sl<23> vdd vss wl<90> / cell_PIM2
XI20004 bl<21> cbl<10> in1<53> in2<53> sl<21> vdd vss wl<53> / cell_PIM2
XI20583 bl<31> cbl<15> in1<21> in2<21> sl<31> vdd vss wl<21> / cell_PIM2
XI19407 bl<23> cbl<11> in1<92> in2<92> sl<23> vdd vss wl<92> / cell_PIM2
XI19406 bl<23> cbl<11> in1<93> in2<93> sl<23> vdd vss wl<93> / cell_PIM2
XI19408 bl<23> cbl<11> in1<91> in2<91> sl<23> vdd vss wl<91> / cell_PIM2
XI19998 bl<19> cbl<9> in1<51> in2<51> sl<19> vdd vss wl<51> / cell_PIM2
XI19997 bl<19> cbl<9> in1<52> in2<52> sl<19> vdd vss wl<52> / cell_PIM2
XI20578 bl<29> cbl<14> in1<19> in2<19> sl<29> vdd vss wl<19> / cell_PIM2
XI20577 bl<29> cbl<14> in1<18> in2<18> sl<29> vdd vss wl<18> / cell_PIM2
XI20576 bl<29> cbl<14> in1<21> in2<21> sl<29> vdd vss wl<21> / cell_PIM2
XI20575 bl<29> cbl<14> in1<20> in2<20> sl<29> vdd vss wl<20> / cell_PIM2
XI19400 bl<21> cbl<10> in1<91> in2<91> sl<21> vdd vss wl<91> / cell_PIM2
XI19399 bl<21> cbl<10> in1<90> in2<90> sl<21> vdd vss wl<90> / cell_PIM2
XI19996 bl<19> cbl<9> in1<53> in2<53> sl<19> vdd vss wl<53> / cell_PIM2
XI19995 bl<19> cbl<9> in1<54> in2<54> sl<19> vdd vss wl<54> / cell_PIM2
XI19994 bl<19> cbl<9> in1<55> in2<55> sl<19> vdd vss wl<55> / cell_PIM2
XI20570 bl<27> cbl<13> in1<18> in2<18> sl<27> vdd vss wl<18> / cell_PIM2
XI20569 bl<27> cbl<13> in1<19> in2<19> sl<27> vdd vss wl<19> / cell_PIM2
XI20568 bl<27> cbl<13> in1<20> in2<20> sl<27> vdd vss wl<20> / cell_PIM2
XI20567 bl<27> cbl<13> in1<21> in2<21> sl<27> vdd vss wl<21> / cell_PIM2
XI19398 bl<21> cbl<10> in1<89> in2<89> sl<21> vdd vss wl<89> / cell_PIM2
XI19397 bl<21> cbl<10> in1<93> in2<93> sl<21> vdd vss wl<93> / cell_PIM2
XI19396 bl<21> cbl<10> in1<92> in2<92> sl<21> vdd vss wl<92> / cell_PIM2
XI19390 bl<19> cbl<9> in1<89> in2<89> sl<19> vdd vss wl<89> / cell_PIM2
XI19389 bl<19> cbl<9> in1<90> in2<90> sl<19> vdd vss wl<90> / cell_PIM2
XI19988 bl<17> cbl<8> in1<52> in2<52> sl<17> vdd vss wl<52> / cell_PIM2
XI19987 bl<17> cbl<8> in1<51> in2<51> sl<17> vdd vss wl<51> / cell_PIM2
XI19986 bl<17> cbl<8> in1<55> in2<55> sl<17> vdd vss wl<55> / cell_PIM2
XI19985 bl<17> cbl<8> in1<54> in2<54> sl<17> vdd vss wl<54> / cell_PIM2
XI20562 bl<25> cbl<12> in1<18> in2<18> sl<25> vdd vss wl<18> / cell_PIM2
XI20561 bl<25> cbl<12> in1<19> in2<19> sl<25> vdd vss wl<19> / cell_PIM2
XI20560 bl<25> cbl<12> in1<20> in2<20> sl<25> vdd vss wl<20> / cell_PIM2
XI20559 bl<25> cbl<12> in1<21> in2<21> sl<25> vdd vss wl<21> / cell_PIM2
XI19387 bl<19> cbl<9> in1<92> in2<92> sl<19> vdd vss wl<92> / cell_PIM2
XI19386 bl<19> cbl<9> in1<93> in2<93> sl<19> vdd vss wl<93> / cell_PIM2
XI19388 bl<19> cbl<9> in1<91> in2<91> sl<19> vdd vss wl<91> / cell_PIM2
XI19984 bl<17> cbl<8> in1<53> in2<53> sl<17> vdd vss wl<53> / cell_PIM2
XI20554 bl<23> cbl<11> in1<18> in2<18> sl<23> vdd vss wl<18> / cell_PIM2
XI19380 bl<17> cbl<8> in1<91> in2<91> sl<17> vdd vss wl<91> / cell_PIM2
XI19379 bl<17> cbl<8> in1<90> in2<90> sl<17> vdd vss wl<90> / cell_PIM2
XI19978 bl<31> cbl<15> in1<56> in2<56> sl<31> vdd vss wl<56> / cell_PIM2
XI19977 bl<31> cbl<15> in1<57> in2<57> sl<31> vdd vss wl<57> / cell_PIM2
XI20553 bl<23> cbl<11> in1<19> in2<19> sl<23> vdd vss wl<19> / cell_PIM2
XI20552 bl<23> cbl<11> in1<20> in2<20> sl<23> vdd vss wl<20> / cell_PIM2
XI20551 bl<23> cbl<11> in1<21> in2<21> sl<23> vdd vss wl<21> / cell_PIM2
XI20546 bl<21> cbl<10> in1<19> in2<19> sl<21> vdd vss wl<19> / cell_PIM2
XI20545 bl<21> cbl<10> in1<18> in2<18> sl<21> vdd vss wl<18> / cell_PIM2
XI20544 bl<21> cbl<10> in1<21> in2<21> sl<21> vdd vss wl<21> / cell_PIM2
XI19976 bl<31> cbl<15> in1<58> in2<58> sl<31> vdd vss wl<58> / cell_PIM2
XI19975 bl<31> cbl<15> in1<59> in2<59> sl<31> vdd vss wl<59> / cell_PIM2
XI19974 bl<31> cbl<15> in1<60> in2<60> sl<31> vdd vss wl<60> / cell_PIM2
XI19378 bl<17> cbl<8> in1<89> in2<89> sl<17> vdd vss wl<89> / cell_PIM2
XI19377 bl<17> cbl<8> in1<93> in2<93> sl<17> vdd vss wl<93> / cell_PIM2
XI19376 bl<17> cbl<8> in1<92> in2<92> sl<17> vdd vss wl<92> / cell_PIM2
XI19370 bl<31> cbl<15> in1<94> in2<94> sl<31> vdd vss wl<94> / cell_PIM2
XI19369 bl<31> cbl<15> in1<95> in2<95> sl<31> vdd vss wl<95> / cell_PIM2
XI20543 bl<21> cbl<10> in1<20> in2<20> sl<21> vdd vss wl<20> / cell_PIM2
XI19367 bl<31> cbl<15> in1<97> in2<97> sl<31> vdd vss wl<97> / cell_PIM2
XI19366 bl<31> cbl<15> in1<98> in2<98> sl<31> vdd vss wl<98> / cell_PIM2
XI19368 bl<31> cbl<15> in1<96> in2<96> sl<31> vdd vss wl<96> / cell_PIM2
XI19968 bl<29> cbl<14> in1<57> in2<57> sl<29> vdd vss wl<57> / cell_PIM2
XI19967 bl<29> cbl<14> in1<56> in2<56> sl<29> vdd vss wl<56> / cell_PIM2
XI19966 bl<29> cbl<14> in1<60> in2<60> sl<29> vdd vss wl<60> / cell_PIM2
XI19965 bl<29> cbl<14> in1<59> in2<59> sl<29> vdd vss wl<59> / cell_PIM2
XI20538 bl<19> cbl<9> in1<18> in2<18> sl<19> vdd vss wl<18> / cell_PIM2
XI20537 bl<19> cbl<9> in1<19> in2<19> sl<19> vdd vss wl<19> / cell_PIM2
XI20536 bl<19> cbl<9> in1<20> in2<20> sl<19> vdd vss wl<20> / cell_PIM2
XI20535 bl<19> cbl<9> in1<21> in2<21> sl<19> vdd vss wl<21> / cell_PIM2
XI19360 bl<29> cbl<14> in1<95> in2<95> sl<29> vdd vss wl<95> / cell_PIM2
XI19359 bl<29> cbl<14> in1<94> in2<94> sl<29> vdd vss wl<94> / cell_PIM2
XI19964 bl<29> cbl<14> in1<58> in2<58> sl<29> vdd vss wl<58> / cell_PIM2
XI20530 bl<17> cbl<8> in1<19> in2<19> sl<17> vdd vss wl<19> / cell_PIM2
XI20529 bl<17> cbl<8> in1<18> in2<18> sl<17> vdd vss wl<18> / cell_PIM2
XI20528 bl<17> cbl<8> in1<21> in2<21> sl<17> vdd vss wl<21> / cell_PIM2
XI20527 bl<17> cbl<8> in1<20> in2<20> sl<17> vdd vss wl<20> / cell_PIM2
XI19958 bl<27> cbl<13> in1<56> in2<56> sl<27> vdd vss wl<56> / cell_PIM2
XI19957 bl<27> cbl<13> in1<57> in2<57> sl<27> vdd vss wl<57> / cell_PIM2
XI19358 bl<29> cbl<14> in1<98> in2<98> sl<29> vdd vss wl<98> / cell_PIM2
XI19357 bl<29> cbl<14> in1<97> in2<97> sl<29> vdd vss wl<97> / cell_PIM2
XI19356 bl<29> cbl<14> in1<96> in2<96> sl<29> vdd vss wl<96> / cell_PIM2
XI19350 bl<27> cbl<13> in1<94> in2<94> sl<27> vdd vss wl<94> / cell_PIM2
XI19349 bl<27> cbl<13> in1<95> in2<95> sl<27> vdd vss wl<95> / cell_PIM2
XI19956 bl<27> cbl<13> in1<58> in2<58> sl<27> vdd vss wl<58> / cell_PIM2
XI19955 bl<27> cbl<13> in1<59> in2<59> sl<27> vdd vss wl<59> / cell_PIM2
XI19954 bl<27> cbl<13> in1<60> in2<60> sl<27> vdd vss wl<60> / cell_PIM2
XI20522 bl<31> cbl<15> in1<22> in2<22> sl<31> vdd vss wl<22> / cell_PIM2
XI20521 bl<31> cbl<15> in1<23> in2<23> sl<31> vdd vss wl<23> / cell_PIM2
XI20520 bl<31> cbl<15> in1<24> in2<24> sl<31> vdd vss wl<24> / cell_PIM2
XI20519 bl<31> cbl<15> in1<25> in2<25> sl<31> vdd vss wl<25> / cell_PIM2
XI19347 bl<27> cbl<13> in1<97> in2<97> sl<27> vdd vss wl<97> / cell_PIM2
XI19346 bl<27> cbl<13> in1<98> in2<98> sl<27> vdd vss wl<98> / cell_PIM2
XI19348 bl<27> cbl<13> in1<96> in2<96> sl<27> vdd vss wl<96> / cell_PIM2
XI20518 bl<31> cbl<15> in1<26> in2<26> sl<31> vdd vss wl<26> / cell_PIM2
XI19340 bl<25> cbl<12> in1<94> in2<94> sl<25> vdd vss wl<94> / cell_PIM2
XI19339 bl<25> cbl<12> in1<95> in2<95> sl<25> vdd vss wl<95> / cell_PIM2
XI19948 bl<25> cbl<12> in1<56> in2<56> sl<25> vdd vss wl<56> / cell_PIM2
XI19947 bl<25> cbl<12> in1<57> in2<57> sl<25> vdd vss wl<57> / cell_PIM2
XI19946 bl<25> cbl<12> in1<58> in2<58> sl<25> vdd vss wl<58> / cell_PIM2
XI19945 bl<25> cbl<12> in1<59> in2<59> sl<25> vdd vss wl<59> / cell_PIM2
XI20512 bl<29> cbl<14> in1<24> in2<24> sl<29> vdd vss wl<24> / cell_PIM2
XI20511 bl<29> cbl<14> in1<23> in2<23> sl<29> vdd vss wl<23> / cell_PIM2
XI20510 bl<29> cbl<14> in1<22> in2<22> sl<29> vdd vss wl<22> / cell_PIM2
XI20509 bl<29> cbl<14> in1<26> in2<26> sl<29> vdd vss wl<26> / cell_PIM2
XI20508 bl<29> cbl<14> in1<25> in2<25> sl<29> vdd vss wl<25> / cell_PIM2
XI19944 bl<25> cbl<12> in1<60> in2<60> sl<25> vdd vss wl<60> / cell_PIM2
XI19338 bl<25> cbl<12> in1<96> in2<96> sl<25> vdd vss wl<96> / cell_PIM2
XI19337 bl<25> cbl<12> in1<97> in2<97> sl<25> vdd vss wl<97> / cell_PIM2
XI19336 bl<25> cbl<12> in1<98> in2<98> sl<25> vdd vss wl<98> / cell_PIM2
XI19330 bl<23> cbl<11> in1<94> in2<94> sl<23> vdd vss wl<94> / cell_PIM2
XI19329 bl<23> cbl<11> in1<95> in2<95> sl<23> vdd vss wl<95> / cell_PIM2
XI19938 bl<23> cbl<11> in1<56> in2<56> sl<23> vdd vss wl<56> / cell_PIM2
XI19937 bl<23> cbl<11> in1<57> in2<57> sl<23> vdd vss wl<57> / cell_PIM2
XI20502 bl<27> cbl<13> in1<22> in2<22> sl<27> vdd vss wl<22> / cell_PIM2
XI20501 bl<27> cbl<13> in1<23> in2<23> sl<27> vdd vss wl<23> / cell_PIM2
XI20500 bl<27> cbl<13> in1<24> in2<24> sl<27> vdd vss wl<24> / cell_PIM2
XI20499 bl<27> cbl<13> in1<25> in2<25> sl<27> vdd vss wl<25> / cell_PIM2
XI19327 bl<23> cbl<11> in1<97> in2<97> sl<23> vdd vss wl<97> / cell_PIM2
XI19326 bl<23> cbl<11> in1<98> in2<98> sl<23> vdd vss wl<98> / cell_PIM2
XI19328 bl<23> cbl<11> in1<96> in2<96> sl<23> vdd vss wl<96> / cell_PIM2
XI19936 bl<23> cbl<11> in1<58> in2<58> sl<23> vdd vss wl<58> / cell_PIM2
XI19935 bl<23> cbl<11> in1<59> in2<59> sl<23> vdd vss wl<59> / cell_PIM2
XI19934 bl<23> cbl<11> in1<60> in2<60> sl<23> vdd vss wl<60> / cell_PIM2
XI20498 bl<27> cbl<13> in1<26> in2<26> sl<27> vdd vss wl<26> / cell_PIM2
XI19320 bl<21> cbl<10> in1<95> in2<95> sl<21> vdd vss wl<95> / cell_PIM2
XI19319 bl<21> cbl<10> in1<94> in2<94> sl<21> vdd vss wl<94> / cell_PIM2
XI20492 bl<25> cbl<12> in1<22> in2<22> sl<25> vdd vss wl<22> / cell_PIM2
XI20491 bl<25> cbl<12> in1<23> in2<23> sl<25> vdd vss wl<23> / cell_PIM2
XI20490 bl<25> cbl<12> in1<24> in2<24> sl<25> vdd vss wl<24> / cell_PIM2
XI20489 bl<25> cbl<12> in1<25> in2<25> sl<25> vdd vss wl<25> / cell_PIM2
XI20488 bl<25> cbl<12> in1<26> in2<26> sl<25> vdd vss wl<26> / cell_PIM2
XI19928 bl<21> cbl<10> in1<57> in2<57> sl<21> vdd vss wl<57> / cell_PIM2
XI19927 bl<21> cbl<10> in1<56> in2<56> sl<21> vdd vss wl<56> / cell_PIM2
XI19926 bl<21> cbl<10> in1<60> in2<60> sl<21> vdd vss wl<60> / cell_PIM2
XI19925 bl<21> cbl<10> in1<59> in2<59> sl<21> vdd vss wl<59> / cell_PIM2
XI19318 bl<21> cbl<10> in1<98> in2<98> sl<21> vdd vss wl<98> / cell_PIM2
XI19317 bl<21> cbl<10> in1<97> in2<97> sl<21> vdd vss wl<97> / cell_PIM2
XI19316 bl<21> cbl<10> in1<96> in2<96> sl<21> vdd vss wl<96> / cell_PIM2
XI19310 bl<19> cbl<9> in1<94> in2<94> sl<19> vdd vss wl<94> / cell_PIM2
XI19309 bl<19> cbl<9> in1<95> in2<95> sl<19> vdd vss wl<95> / cell_PIM2
XI19924 bl<21> cbl<10> in1<58> in2<58> sl<21> vdd vss wl<58> / cell_PIM2
XI20482 bl<23> cbl<11> in1<22> in2<22> sl<23> vdd vss wl<22> / cell_PIM2
XI20481 bl<23> cbl<11> in1<23> in2<23> sl<23> vdd vss wl<23> / cell_PIM2
XI20480 bl<23> cbl<11> in1<24> in2<24> sl<23> vdd vss wl<24> / cell_PIM2
XI20479 bl<23> cbl<11> in1<25> in2<25> sl<23> vdd vss wl<25> / cell_PIM2
XI19307 bl<19> cbl<9> in1<97> in2<97> sl<19> vdd vss wl<97> / cell_PIM2
XI19306 bl<19> cbl<9> in1<98> in2<98> sl<19> vdd vss wl<98> / cell_PIM2
XI19308 bl<19> cbl<9> in1<96> in2<96> sl<19> vdd vss wl<96> / cell_PIM2
XI19918 bl<19> cbl<9> in1<56> in2<56> sl<19> vdd vss wl<56> / cell_PIM2
XI19917 bl<19> cbl<9> in1<57> in2<57> sl<19> vdd vss wl<57> / cell_PIM2
XI20478 bl<23> cbl<11> in1<26> in2<26> sl<23> vdd vss wl<26> / cell_PIM2
XI19300 bl<17> cbl<8> in1<95> in2<95> sl<17> vdd vss wl<95> / cell_PIM2
XI19299 bl<17> cbl<8> in1<94> in2<94> sl<17> vdd vss wl<94> / cell_PIM2
XI19916 bl<19> cbl<9> in1<58> in2<58> sl<19> vdd vss wl<58> / cell_PIM2
XI19915 bl<19> cbl<9> in1<59> in2<59> sl<19> vdd vss wl<59> / cell_PIM2
XI19914 bl<19> cbl<9> in1<60> in2<60> sl<19> vdd vss wl<60> / cell_PIM2
XI20472 bl<21> cbl<10> in1<24> in2<24> sl<21> vdd vss wl<24> / cell_PIM2
XI20471 bl<21> cbl<10> in1<23> in2<23> sl<21> vdd vss wl<23> / cell_PIM2
XI20470 bl<21> cbl<10> in1<22> in2<22> sl<21> vdd vss wl<22> / cell_PIM2
XI20469 bl<21> cbl<10> in1<26> in2<26> sl<21> vdd vss wl<26> / cell_PIM2
XI20468 bl<21> cbl<10> in1<25> in2<25> sl<21> vdd vss wl<25> / cell_PIM2
XI19298 bl<17> cbl<8> in1<98> in2<98> sl<17> vdd vss wl<98> / cell_PIM2
XI19297 bl<17> cbl<8> in1<97> in2<97> sl<17> vdd vss wl<97> / cell_PIM2
XI19296 bl<17> cbl<8> in1<96> in2<96> sl<17> vdd vss wl<96> / cell_PIM2
XI19290 bl<31> cbl<15> in1<99> in2<99> sl<31> vdd vss wl<99> / cell_PIM2
XI19289 bl<31> cbl<15> in1<100> in2<100> sl<31> vdd vss wl<100> / cell_PIM2
XI19908 bl<17> cbl<8> in1<57> in2<57> sl<17> vdd vss wl<57> / cell_PIM2
XI19907 bl<17> cbl<8> in1<56> in2<56> sl<17> vdd vss wl<56> / cell_PIM2
XI19906 bl<17> cbl<8> in1<60> in2<60> sl<17> vdd vss wl<60> / cell_PIM2
XI19905 bl<17> cbl<8> in1<59> in2<59> sl<17> vdd vss wl<59> / cell_PIM2
XI20462 bl<19> cbl<9> in1<22> in2<22> sl<19> vdd vss wl<22> / cell_PIM2
XI20461 bl<19> cbl<9> in1<23> in2<23> sl<19> vdd vss wl<23> / cell_PIM2
XI20460 bl<19> cbl<9> in1<24> in2<24> sl<19> vdd vss wl<24> / cell_PIM2
XI20459 bl<19> cbl<9> in1<25> in2<25> sl<19> vdd vss wl<25> / cell_PIM2
XI19287 bl<31> cbl<15> in1<102> in2<102> sl<31> vdd vss wl<102> / cell_PIM2
XI19286 bl<31> cbl<15> in1<103> in2<103> sl<31> vdd vss wl<103> / cell_PIM2
XI19288 bl<31> cbl<15> in1<101> in2<101> sl<31> vdd vss wl<101> / cell_PIM2
XI19904 bl<17> cbl<8> in1<58> in2<58> sl<17> vdd vss wl<58> / cell_PIM2
XI20458 bl<19> cbl<9> in1<26> in2<26> sl<19> vdd vss wl<26> / cell_PIM2
XI17493 bl<7> cbl<3> in1<78> in2<78> sl<7> vdd vss wl<78> / cell_PIM2
XI17492 bl<7> cbl<3> in1<79> in2<79> sl<7> vdd vss wl<79> / cell_PIM2
XI17491 bl<7> cbl<3> in1<80> in2<80> sl<7> vdd vss wl<80> / cell_PIM2
XI17490 bl<7> cbl<3> in1<81> in2<81> sl<7> vdd vss wl<81> / cell_PIM2
XI18140 bl<9> cbl<4> in1<86> in2<86> sl<9> vdd vss wl<86> / cell_PIM2
XI18139 bl<9> cbl<4> in1<85> in2<85> sl<9> vdd vss wl<85> / cell_PIM2
XI18793 bl<9> cbl<4> in1<3> in2<3> sl<9> vdd vss wl<3> / cell_PIM2
XI18792 bl<9> cbl<4> in1<4> in2<4> sl<9> vdd vss wl<4> / cell_PIM2
XI18791 bl<9> cbl<4> in1<1> in2<1> sl<9> vdd vss wl<1> / cell_PIM2
XI18786 bl<15> cbl<7> in1<5> in2<5> sl<15> vdd vss wl<5> / cell_PIM2
XI18785 bl<15> cbl<7> in1<6> in2<6> sl<15> vdd vss wl<6> / cell_PIM2
XI18784 bl<15> cbl<7> in1<7> in2<7> sl<15> vdd vss wl<7> / cell_PIM2
XI18138 bl<9> cbl<4> in1<84> in2<84> sl<9> vdd vss wl<84> / cell_PIM2
XI18137 bl<9> cbl<4> in1<83> in2<83> sl<9> vdd vss wl<83> / cell_PIM2
XI18136 bl<9> cbl<4> in1<82> in2<82> sl<9> vdd vss wl<82> / cell_PIM2
XI17484 bl<5> cbl<2> in1<81> in2<81> sl<5> vdd vss wl<81> / cell_PIM2
XI17483 bl<5> cbl<2> in1<80> in2<80> sl<5> vdd vss wl<80> / cell_PIM2
XI17482 bl<5> cbl<2> in1<79> in2<79> sl<5> vdd vss wl<79> / cell_PIM2
XI17481 bl<5> cbl<2> in1<78> in2<78> sl<5> vdd vss wl<78> / cell_PIM2
XI17480 bl<5> cbl<2> in1<77> in2<77> sl<5> vdd vss wl<77> / cell_PIM2
XI18130 bl<15> cbl<7> in1<87> in2<87> sl<15> vdd vss wl<87> / cell_PIM2
XI18129 bl<15> cbl<7> in1<88> in2<88> sl<15> vdd vss wl<88> / cell_PIM2
XI18783 bl<15> cbl<7> in1<8> in2<8> sl<15> vdd vss wl<8> / cell_PIM2
XI18782 bl<15> cbl<7> in1<9> in2<9> sl<15> vdd vss wl<9> / cell_PIM2
XI17474 bl<7> cbl<3> in1<82> in2<82> sl<7> vdd vss wl<82> / cell_PIM2
XI18128 bl<15> cbl<7> in1<89> in2<89> sl<15> vdd vss wl<89> / cell_PIM2
XI18127 bl<15> cbl<7> in1<90> in2<90> sl<15> vdd vss wl<90> / cell_PIM2
XI18126 bl<15> cbl<7> in1<91> in2<91> sl<15> vdd vss wl<91> / cell_PIM2
XI18776 bl<13> cbl<6> in1<9> in2<9> sl<13> vdd vss wl<9> / cell_PIM2
XI18775 bl<13> cbl<6> in1<8> in2<8> sl<13> vdd vss wl<8> / cell_PIM2
XI18774 bl<13> cbl<6> in1<7> in2<7> sl<13> vdd vss wl<7> / cell_PIM2
XI17473 bl<7> cbl<3> in1<83> in2<83> sl<7> vdd vss wl<83> / cell_PIM2
XI17472 bl<7> cbl<3> in1<84> in2<84> sl<7> vdd vss wl<84> / cell_PIM2
XI17471 bl<7> cbl<3> in1<85> in2<85> sl<7> vdd vss wl<85> / cell_PIM2
XI17470 bl<7> cbl<3> in1<86> in2<86> sl<7> vdd vss wl<86> / cell_PIM2
XI18120 bl<13> cbl<6> in1<91> in2<91> sl<13> vdd vss wl<91> / cell_PIM2
XI18119 bl<13> cbl<6> in1<90> in2<90> sl<13> vdd vss wl<90> / cell_PIM2
XI18773 bl<13> cbl<6> in1<6> in2<6> sl<13> vdd vss wl<6> / cell_PIM2
XI18772 bl<13> cbl<6> in1<5> in2<5> sl<13> vdd vss wl<5> / cell_PIM2
XI18766 bl<11> cbl<5> in1<5> in2<5> sl<11> vdd vss wl<5> / cell_PIM2
XI18765 bl<11> cbl<5> in1<6> in2<6> sl<11> vdd vss wl<6> / cell_PIM2
XI18764 bl<11> cbl<5> in1<7> in2<7> sl<11> vdd vss wl<7> / cell_PIM2
XI18118 bl<13> cbl<6> in1<89> in2<89> sl<13> vdd vss wl<89> / cell_PIM2
XI18117 bl<13> cbl<6> in1<88> in2<88> sl<13> vdd vss wl<88> / cell_PIM2
XI18116 bl<13> cbl<6> in1<87> in2<87> sl<13> vdd vss wl<87> / cell_PIM2
XI17464 bl<5> cbl<2> in1<86> in2<86> sl<5> vdd vss wl<86> / cell_PIM2
XI17463 bl<5> cbl<2> in1<85> in2<85> sl<5> vdd vss wl<85> / cell_PIM2
XI17462 bl<5> cbl<2> in1<84> in2<84> sl<5> vdd vss wl<84> / cell_PIM2
XI17461 bl<5> cbl<2> in1<83> in2<83> sl<5> vdd vss wl<83> / cell_PIM2
XI17460 bl<5> cbl<2> in1<82> in2<82> sl<5> vdd vss wl<82> / cell_PIM2
XI18110 bl<11> cbl<5> in1<87> in2<87> sl<11> vdd vss wl<87> / cell_PIM2
XI18109 bl<11> cbl<5> in1<88> in2<88> sl<11> vdd vss wl<88> / cell_PIM2
XI18763 bl<11> cbl<5> in1<8> in2<8> sl<11> vdd vss wl<8> / cell_PIM2
XI18762 bl<11> cbl<5> in1<9> in2<9> sl<11> vdd vss wl<9> / cell_PIM2
XI17454 bl<7> cbl<3> in1<87> in2<87> sl<7> vdd vss wl<87> / cell_PIM2
XI18108 bl<11> cbl<5> in1<89> in2<89> sl<11> vdd vss wl<89> / cell_PIM2
XI18107 bl<11> cbl<5> in1<90> in2<90> sl<11> vdd vss wl<90> / cell_PIM2
XI18106 bl<11> cbl<5> in1<91> in2<91> sl<11> vdd vss wl<91> / cell_PIM2
XI18756 bl<9> cbl<4> in1<9> in2<9> sl<9> vdd vss wl<9> / cell_PIM2
XI18755 bl<9> cbl<4> in1<8> in2<8> sl<9> vdd vss wl<8> / cell_PIM2
XI18754 bl<9> cbl<4> in1<7> in2<7> sl<9> vdd vss wl<7> / cell_PIM2
XI17453 bl<7> cbl<3> in1<88> in2<88> sl<7> vdd vss wl<88> / cell_PIM2
XI17452 bl<7> cbl<3> in1<89> in2<89> sl<7> vdd vss wl<89> / cell_PIM2
XI17451 bl<7> cbl<3> in1<90> in2<90> sl<7> vdd vss wl<90> / cell_PIM2
XI17450 bl<7> cbl<3> in1<91> in2<91> sl<7> vdd vss wl<91> / cell_PIM2
XI18100 bl<9> cbl<4> in1<91> in2<91> sl<9> vdd vss wl<91> / cell_PIM2
XI18099 bl<9> cbl<4> in1<90> in2<90> sl<9> vdd vss wl<90> / cell_PIM2
XI18753 bl<9> cbl<4> in1<6> in2<6> sl<9> vdd vss wl<6> / cell_PIM2
XI18752 bl<9> cbl<4> in1<5> in2<5> sl<9> vdd vss wl<5> / cell_PIM2
XI18746 bl<15> cbl<7> in1<10> in2<10> sl<15> vdd vss wl<10> / cell_PIM2
XI18745 bl<15> cbl<7> in1<11> in2<11> sl<15> vdd vss wl<11> / cell_PIM2
XI18744 bl<15> cbl<7> in1<12> in2<12> sl<15> vdd vss wl<12> / cell_PIM2
XI18098 bl<9> cbl<4> in1<89> in2<89> sl<9> vdd vss wl<89> / cell_PIM2
XI18097 bl<9> cbl<4> in1<88> in2<88> sl<9> vdd vss wl<88> / cell_PIM2
XI18096 bl<9> cbl<4> in1<87> in2<87> sl<9> vdd vss wl<87> / cell_PIM2
XI17444 bl<5> cbl<2> in1<91> in2<91> sl<5> vdd vss wl<91> / cell_PIM2
XI17443 bl<5> cbl<2> in1<90> in2<90> sl<5> vdd vss wl<90> / cell_PIM2
XI17442 bl<5> cbl<2> in1<89> in2<89> sl<5> vdd vss wl<89> / cell_PIM2
XI17441 bl<5> cbl<2> in1<88> in2<88> sl<5> vdd vss wl<88> / cell_PIM2
XI17440 bl<5> cbl<2> in1<87> in2<87> sl<5> vdd vss wl<87> / cell_PIM2
XI18090 bl<15> cbl<7> in1<92> in2<92> sl<15> vdd vss wl<92> / cell_PIM2
XI18089 bl<15> cbl<7> in1<93> in2<93> sl<15> vdd vss wl<93> / cell_PIM2
XI18743 bl<15> cbl<7> in1<13> in2<13> sl<15> vdd vss wl<13> / cell_PIM2
XI18742 bl<15> cbl<7> in1<14> in2<14> sl<15> vdd vss wl<14> / cell_PIM2
XI17434 bl<7> cbl<3> in1<92> in2<92> sl<7> vdd vss wl<92> / cell_PIM2
XI18088 bl<15> cbl<7> in1<94> in2<94> sl<15> vdd vss wl<94> / cell_PIM2
XI18087 bl<15> cbl<7> in1<95> in2<95> sl<15> vdd vss wl<95> / cell_PIM2
XI18736 bl<13> cbl<6> in1<14> in2<14> sl<13> vdd vss wl<14> / cell_PIM2
XI18735 bl<13> cbl<6> in1<13> in2<13> sl<13> vdd vss wl<13> / cell_PIM2
XI18734 bl<13> cbl<6> in1<12> in2<12> sl<13> vdd vss wl<12> / cell_PIM2
XI17433 bl<7> cbl<3> in1<93> in2<93> sl<7> vdd vss wl<93> / cell_PIM2
XI17432 bl<7> cbl<3> in1<94> in2<94> sl<7> vdd vss wl<94> / cell_PIM2
XI17431 bl<7> cbl<3> in1<95> in2<95> sl<7> vdd vss wl<95> / cell_PIM2
XI18082 bl<13> cbl<6> in1<95> in2<95> sl<13> vdd vss wl<95> / cell_PIM2
XI18081 bl<13> cbl<6> in1<94> in2<94> sl<13> vdd vss wl<94> / cell_PIM2
XI18080 bl<13> cbl<6> in1<93> in2<93> sl<13> vdd vss wl<93> / cell_PIM2
XI18079 bl<13> cbl<6> in1<92> in2<92> sl<13> vdd vss wl<92> / cell_PIM2
XI18733 bl<13> cbl<6> in1<11> in2<11> sl<13> vdd vss wl<11> / cell_PIM2
XI18732 bl<13> cbl<6> in1<10> in2<10> sl<13> vdd vss wl<10> / cell_PIM2
XI18726 bl<11> cbl<5> in1<10> in2<10> sl<11> vdd vss wl<10> / cell_PIM2
XI18725 bl<11> cbl<5> in1<11> in2<11> sl<11> vdd vss wl<11> / cell_PIM2
XI18724 bl<11> cbl<5> in1<12> in2<12> sl<11> vdd vss wl<12> / cell_PIM2
XI18074 bl<11> cbl<5> in1<92> in2<92> sl<11> vdd vss wl<92> / cell_PIM2
XI17426 bl<5> cbl<2> in1<95> in2<95> sl<5> vdd vss wl<95> / cell_PIM2
XI17425 bl<5> cbl<2> in1<94> in2<94> sl<5> vdd vss wl<94> / cell_PIM2
XI17424 bl<5> cbl<2> in1<93> in2<93> sl<5> vdd vss wl<93> / cell_PIM2
XI17423 bl<5> cbl<2> in1<92> in2<92> sl<5> vdd vss wl<92> / cell_PIM2
XI18073 bl<11> cbl<5> in1<93> in2<93> sl<11> vdd vss wl<93> / cell_PIM2
XI18072 bl<11> cbl<5> in1<94> in2<94> sl<11> vdd vss wl<94> / cell_PIM2
XI18071 bl<11> cbl<5> in1<95> in2<95> sl<11> vdd vss wl<95> / cell_PIM2
XI18723 bl<11> cbl<5> in1<13> in2<13> sl<11> vdd vss wl<13> / cell_PIM2
XI18722 bl<11> cbl<5> in1<14> in2<14> sl<11> vdd vss wl<14> / cell_PIM2
XI17418 bl<7> cbl<3> in1<96> in2<96> sl<7> vdd vss wl<96> / cell_PIM2
XI17417 bl<7> cbl<3> in1<97> in2<97> sl<7> vdd vss wl<97> / cell_PIM2
XI17416 bl<7> cbl<3> in1<98> in2<98> sl<7> vdd vss wl<98> / cell_PIM2
XI17415 bl<7> cbl<3> in1<99> in2<99> sl<7> vdd vss wl<99> / cell_PIM2
XI17414 bl<7> cbl<3> in1<100> in2<100> sl<7> vdd vss wl<100> / cell_PIM2
XI18066 bl<9> cbl<4> in1<95> in2<95> sl<9> vdd vss wl<95> / cell_PIM2
XI18065 bl<9> cbl<4> in1<94> in2<94> sl<9> vdd vss wl<94> / cell_PIM2
XI18064 bl<9> cbl<4> in1<93> in2<93> sl<9> vdd vss wl<93> / cell_PIM2
XI18716 bl<9> cbl<4> in1<14> in2<14> sl<9> vdd vss wl<14> / cell_PIM2
XI18715 bl<9> cbl<4> in1<13> in2<13> sl<9> vdd vss wl<13> / cell_PIM2
XI18714 bl<9> cbl<4> in1<12> in2<12> sl<9> vdd vss wl<12> / cell_PIM2
XI18063 bl<9> cbl<4> in1<92> in2<92> sl<9> vdd vss wl<92> / cell_PIM2
XI18713 bl<9> cbl<4> in1<11> in2<11> sl<9> vdd vss wl<11> / cell_PIM2
XI18712 bl<9> cbl<4> in1<10> in2<10> sl<9> vdd vss wl<10> / cell_PIM2
XI18706 bl<15> cbl<7> in1<15> in2<15> sl<15> vdd vss wl<15> / cell_PIM2
XI18705 bl<15> cbl<7> in1<16> in2<16> sl<15> vdd vss wl<16> / cell_PIM2
XI18704 bl<15> cbl<7> in1<17> in2<17> sl<15> vdd vss wl<17> / cell_PIM2
XI18058 bl<15> cbl<7> in1<96> in2<96> sl<15> vdd vss wl<96> / cell_PIM2
XI18057 bl<15> cbl<7> in1<97> in2<97> sl<15> vdd vss wl<97> / cell_PIM2
XI18056 bl<15> cbl<7> in1<98> in2<98> sl<15> vdd vss wl<98> / cell_PIM2
XI18055 bl<15> cbl<7> in1<99> in2<99> sl<15> vdd vss wl<99> / cell_PIM2
XI18054 bl<15> cbl<7> in1<100> in2<100> sl<15> vdd vss wl<100> / cell_PIM2
XI17408 bl<5> cbl<2> in1<100> in2<100> sl<5> vdd vss wl<100> / cell_PIM2
XI17407 bl<5> cbl<2> in1<99> in2<99> sl<5> vdd vss wl<99> / cell_PIM2
XI17406 bl<5> cbl<2> in1<98> in2<98> sl<5> vdd vss wl<98> / cell_PIM2
XI17405 bl<5> cbl<2> in1<97> in2<97> sl<5> vdd vss wl<97> / cell_PIM2
XI17404 bl<5> cbl<2> in1<96> in2<96> sl<5> vdd vss wl<96> / cell_PIM2
XI18703 bl<15> cbl<7> in1<18> in2<18> sl<15> vdd vss wl<18> / cell_PIM2
XI18702 bl<15> cbl<7> in1<19> in2<19> sl<15> vdd vss wl<19> / cell_PIM2
XI17398 bl<7> cbl<3> in1<101> in2<101> sl<7> vdd vss wl<101> / cell_PIM2
XI17397 bl<7> cbl<3> in1<102> in2<102> sl<7> vdd vss wl<102> / cell_PIM2
XI17396 bl<7> cbl<3> in1<103> in2<103> sl<7> vdd vss wl<103> / cell_PIM2
XI17395 bl<7> cbl<3> in1<104> in2<104> sl<7> vdd vss wl<104> / cell_PIM2
XI17394 bl<7> cbl<3> in1<105> in2<105> sl<7> vdd vss wl<105> / cell_PIM2
XI18048 bl<13> cbl<6> in1<100> in2<100> sl<13> vdd vss wl<100> / cell_PIM2
XI18047 bl<13> cbl<6> in1<99> in2<99> sl<13> vdd vss wl<99> / cell_PIM2
XI18046 bl<13> cbl<6> in1<98> in2<98> sl<13> vdd vss wl<98> / cell_PIM2
XI18045 bl<13> cbl<6> in1<97> in2<97> sl<13> vdd vss wl<97> / cell_PIM2
XI18044 bl<13> cbl<6> in1<96> in2<96> sl<13> vdd vss wl<96> / cell_PIM2
XI18696 bl<13> cbl<6> in1<19> in2<19> sl<13> vdd vss wl<19> / cell_PIM2
XI18695 bl<13> cbl<6> in1<18> in2<18> sl<13> vdd vss wl<18> / cell_PIM2
XI18694 bl<13> cbl<6> in1<17> in2<17> sl<13> vdd vss wl<17> / cell_PIM2
XI18693 bl<13> cbl<6> in1<16> in2<16> sl<13> vdd vss wl<16> / cell_PIM2
XI18692 bl<13> cbl<6> in1<15> in2<15> sl<13> vdd vss wl<15> / cell_PIM2
XI18686 bl<11> cbl<5> in1<15> in2<15> sl<11> vdd vss wl<15> / cell_PIM2
XI18685 bl<11> cbl<5> in1<16> in2<16> sl<11> vdd vss wl<16> / cell_PIM2
XI18684 bl<11> cbl<5> in1<17> in2<17> sl<11> vdd vss wl<17> / cell_PIM2
XI18038 bl<11> cbl<5> in1<96> in2<96> sl<11> vdd vss wl<96> / cell_PIM2
XI18037 bl<11> cbl<5> in1<97> in2<97> sl<11> vdd vss wl<97> / cell_PIM2
XI18036 bl<11> cbl<5> in1<98> in2<98> sl<11> vdd vss wl<98> / cell_PIM2
XI18035 bl<11> cbl<5> in1<99> in2<99> sl<11> vdd vss wl<99> / cell_PIM2
XI18034 bl<11> cbl<5> in1<100> in2<100> sl<11> vdd vss wl<100> / cell_PIM2
XI17388 bl<5> cbl<2> in1<105> in2<105> sl<5> vdd vss wl<105> / cell_PIM2
XI17387 bl<5> cbl<2> in1<104> in2<104> sl<5> vdd vss wl<104> / cell_PIM2
XI17386 bl<5> cbl<2> in1<103> in2<103> sl<5> vdd vss wl<103> / cell_PIM2
XI17385 bl<5> cbl<2> in1<102> in2<102> sl<5> vdd vss wl<102> / cell_PIM2
XI17384 bl<5> cbl<2> in1<101> in2<101> sl<5> vdd vss wl<101> / cell_PIM2
XI18683 bl<11> cbl<5> in1<18> in2<18> sl<11> vdd vss wl<18> / cell_PIM2
XI18682 bl<11> cbl<5> in1<19> in2<19> sl<11> vdd vss wl<19> / cell_PIM2
XI17378 bl<7> cbl<3> in1<106> in2<106> sl<7> vdd vss wl<106> / cell_PIM2
XI17377 bl<7> cbl<3> in1<107> in2<107> sl<7> vdd vss wl<107> / cell_PIM2
XI17376 bl<7> cbl<3> in1<108> in2<108> sl<7> vdd vss wl<108> / cell_PIM2
XI17375 bl<7> cbl<3> in1<109> in2<109> sl<7> vdd vss wl<109> / cell_PIM2
XI17374 bl<7> cbl<3> in1<110> in2<110> sl<7> vdd vss wl<110> / cell_PIM2
XI18028 bl<9> cbl<4> in1<100> in2<100> sl<9> vdd vss wl<100> / cell_PIM2
XI18027 bl<9> cbl<4> in1<99> in2<99> sl<9> vdd vss wl<99> / cell_PIM2
XI18026 bl<9> cbl<4> in1<98> in2<98> sl<9> vdd vss wl<98> / cell_PIM2
XI18025 bl<9> cbl<4> in1<97> in2<97> sl<9> vdd vss wl<97> / cell_PIM2
XI18024 bl<9> cbl<4> in1<96> in2<96> sl<9> vdd vss wl<96> / cell_PIM2
XI18676 bl<9> cbl<4> in1<19> in2<19> sl<9> vdd vss wl<19> / cell_PIM2
XI18675 bl<9> cbl<4> in1<18> in2<18> sl<9> vdd vss wl<18> / cell_PIM2
XI18674 bl<9> cbl<4> in1<17> in2<17> sl<9> vdd vss wl<17> / cell_PIM2
XI18673 bl<9> cbl<4> in1<16> in2<16> sl<9> vdd vss wl<16> / cell_PIM2
XI18672 bl<9> cbl<4> in1<15> in2<15> sl<9> vdd vss wl<15> / cell_PIM2
XI18666 bl<15> cbl<7> in1<20> in2<20> sl<15> vdd vss wl<20> / cell_PIM2
XI18665 bl<15> cbl<7> in1<21> in2<21> sl<15> vdd vss wl<21> / cell_PIM2
XI18664 bl<15> cbl<7> in1<22> in2<22> sl<15> vdd vss wl<22> / cell_PIM2
XI18018 bl<15> cbl<7> in1<101> in2<101> sl<15> vdd vss wl<101> / cell_PIM2
XI18017 bl<15> cbl<7> in1<102> in2<102> sl<15> vdd vss wl<102> / cell_PIM2
XI18016 bl<15> cbl<7> in1<103> in2<103> sl<15> vdd vss wl<103> / cell_PIM2
XI18015 bl<15> cbl<7> in1<104> in2<104> sl<15> vdd vss wl<104> / cell_PIM2
XI18014 bl<15> cbl<7> in1<105> in2<105> sl<15> vdd vss wl<105> / cell_PIM2
XI17368 bl<5> cbl<2> in1<110> in2<110> sl<5> vdd vss wl<110> / cell_PIM2
XI17367 bl<5> cbl<2> in1<109> in2<109> sl<5> vdd vss wl<109> / cell_PIM2
XI17366 bl<5> cbl<2> in1<108> in2<108> sl<5> vdd vss wl<108> / cell_PIM2
XI17365 bl<5> cbl<2> in1<107> in2<107> sl<5> vdd vss wl<107> / cell_PIM2
XI17364 bl<5> cbl<2> in1<106> in2<106> sl<5> vdd vss wl<106> / cell_PIM2
XI18663 bl<15> cbl<7> in1<23> in2<23> sl<15> vdd vss wl<23> / cell_PIM2
XI18662 bl<15> cbl<7> in1<24> in2<24> sl<15> vdd vss wl<24> / cell_PIM2
XI17358 bl<7> cbl<3> in1<111> in2<111> sl<7> vdd vss wl<111> / cell_PIM2
XI17357 bl<7> cbl<3> in1<112> in2<112> sl<7> vdd vss wl<112> / cell_PIM2
XI17356 bl<7> cbl<3> in1<113> in2<113> sl<7> vdd vss wl<113> / cell_PIM2
XI17355 bl<7> cbl<3> in1<114> in2<114> sl<7> vdd vss wl<114> / cell_PIM2
XI17354 bl<7> cbl<3> in1<115> in2<115> sl<7> vdd vss wl<115> / cell_PIM2
XI18008 bl<13> cbl<6> in1<105> in2<105> sl<13> vdd vss wl<105> / cell_PIM2
XI18007 bl<13> cbl<6> in1<104> in2<104> sl<13> vdd vss wl<104> / cell_PIM2
XI18006 bl<13> cbl<6> in1<103> in2<103> sl<13> vdd vss wl<103> / cell_PIM2
XI18005 bl<13> cbl<6> in1<102> in2<102> sl<13> vdd vss wl<102> / cell_PIM2
XI18004 bl<13> cbl<6> in1<101> in2<101> sl<13> vdd vss wl<101> / cell_PIM2
XI18656 bl<13> cbl<6> in1<24> in2<24> sl<13> vdd vss wl<24> / cell_PIM2
XI18655 bl<13> cbl<6> in1<23> in2<23> sl<13> vdd vss wl<23> / cell_PIM2
XI18654 bl<13> cbl<6> in1<22> in2<22> sl<13> vdd vss wl<22> / cell_PIM2
XI18653 bl<13> cbl<6> in1<21> in2<21> sl<13> vdd vss wl<21> / cell_PIM2
XI18652 bl<13> cbl<6> in1<20> in2<20> sl<13> vdd vss wl<20> / cell_PIM2
XI18646 bl<11> cbl<5> in1<20> in2<20> sl<11> vdd vss wl<20> / cell_PIM2
XI18645 bl<11> cbl<5> in1<21> in2<21> sl<11> vdd vss wl<21> / cell_PIM2
XI18644 bl<11> cbl<5> in1<22> in2<22> sl<11> vdd vss wl<22> / cell_PIM2
XI17998 bl<11> cbl<5> in1<101> in2<101> sl<11> vdd vss wl<101> / cell_PIM2
XI17997 bl<11> cbl<5> in1<102> in2<102> sl<11> vdd vss wl<102> / cell_PIM2
XI17996 bl<11> cbl<5> in1<103> in2<103> sl<11> vdd vss wl<103> / cell_PIM2
XI17995 bl<11> cbl<5> in1<104> in2<104> sl<11> vdd vss wl<104> / cell_PIM2
XI17994 bl<11> cbl<5> in1<105> in2<105> sl<11> vdd vss wl<105> / cell_PIM2
XI17348 bl<5> cbl<2> in1<115> in2<115> sl<5> vdd vss wl<115> / cell_PIM2
XI17347 bl<5> cbl<2> in1<114> in2<114> sl<5> vdd vss wl<114> / cell_PIM2
XI17346 bl<5> cbl<2> in1<113> in2<113> sl<5> vdd vss wl<113> / cell_PIM2
XI17345 bl<5> cbl<2> in1<112> in2<112> sl<5> vdd vss wl<112> / cell_PIM2
XI17344 bl<5> cbl<2> in1<111> in2<111> sl<5> vdd vss wl<111> / cell_PIM2
XI18643 bl<11> cbl<5> in1<23> in2<23> sl<11> vdd vss wl<23> / cell_PIM2
XI18642 bl<11> cbl<5> in1<24> in2<24> sl<11> vdd vss wl<24> / cell_PIM2
XI17338 bl<7> cbl<3> in1<116> in2<116> sl<7> vdd vss wl<116> / cell_PIM2
XI17337 bl<7> cbl<3> in1<117> in2<117> sl<7> vdd vss wl<117> / cell_PIM2
XI17336 bl<7> cbl<3> in1<118> in2<118> sl<7> vdd vss wl<118> / cell_PIM2
XI17335 bl<7> cbl<3> in1<119> in2<119> sl<7> vdd vss wl<119> / cell_PIM2
XI17988 bl<9> cbl<4> in1<105> in2<105> sl<9> vdd vss wl<105> / cell_PIM2
XI17987 bl<9> cbl<4> in1<104> in2<104> sl<9> vdd vss wl<104> / cell_PIM2
XI17986 bl<9> cbl<4> in1<103> in2<103> sl<9> vdd vss wl<103> / cell_PIM2
XI17985 bl<9> cbl<4> in1<102> in2<102> sl<9> vdd vss wl<102> / cell_PIM2
XI17984 bl<9> cbl<4> in1<101> in2<101> sl<9> vdd vss wl<101> / cell_PIM2
XI18636 bl<9> cbl<4> in1<24> in2<24> sl<9> vdd vss wl<24> / cell_PIM2
XI18635 bl<9> cbl<4> in1<23> in2<23> sl<9> vdd vss wl<23> / cell_PIM2
XI18634 bl<9> cbl<4> in1<22> in2<22> sl<9> vdd vss wl<22> / cell_PIM2
XI24223 bl<55> cbl<27> in1<25> in2<25> sl<55> vdd vss wl<25> / cell_PIM2
XI24872 bl<63> cbl<31> in1<5> in2<5> sl<63> vdd vss wl<5> / cell_PIM2
XI24871 bl<63> cbl<31> in1<6> in2<6> sl<63> vdd vss wl<6> / cell_PIM2
XI24870 bl<63> cbl<31> in1<7> in2<7> sl<63> vdd vss wl<7> / cell_PIM2
XI24873 bl<63> cbl<31> in1<3> in2<3> sl<63> vdd vss wl<3> / cell_PIM2
XI24864 bl<61> cbl<30> in1<3> in2<3> sl<61> vdd vss wl<3> / cell_PIM2
XI24213 bl<53> cbl<26> in1<26> in2<26> sl<53> vdd vss wl<26> / cell_PIM2
XI24862 bl<61> cbl<30> in1<7> in2<7> sl<61> vdd vss wl<7> / cell_PIM2
XI24861 bl<61> cbl<30> in1<6> in2<6> sl<61> vdd vss wl<6> / cell_PIM2
XI24860 bl<61> cbl<30> in1<5> in2<5> sl<61> vdd vss wl<5> / cell_PIM2
XI24863 bl<61> cbl<30> in1<4> in2<4> sl<61> vdd vss wl<4> / cell_PIM2
XI24854 bl<59> cbl<29> in1<4> in2<4> sl<59> vdd vss wl<4> / cell_PIM2
XI24203 bl<51> cbl<25> in1<25> in2<25> sl<51> vdd vss wl<25> / cell_PIM2
XI24852 bl<59> cbl<29> in1<5> in2<5> sl<59> vdd vss wl<5> / cell_PIM2
XI24851 bl<59> cbl<29> in1<6> in2<6> sl<59> vdd vss wl<6> / cell_PIM2
XI24850 bl<59> cbl<29> in1<7> in2<7> sl<59> vdd vss wl<7> / cell_PIM2
XI24853 bl<59> cbl<29> in1<3> in2<3> sl<59> vdd vss wl<3> / cell_PIM2
XI24844 bl<57> cbl<28> in1<4> in2<4> sl<57> vdd vss wl<4> / cell_PIM2
XI24193 bl<49> cbl<24> in1<26> in2<26> sl<49> vdd vss wl<26> / cell_PIM2
XI24842 bl<57> cbl<28> in1<5> in2<5> sl<57> vdd vss wl<5> / cell_PIM2
XI24841 bl<57> cbl<28> in1<6> in2<6> sl<57> vdd vss wl<6> / cell_PIM2
XI24840 bl<57> cbl<28> in1<7> in2<7> sl<57> vdd vss wl<7> / cell_PIM2
XI24843 bl<57> cbl<28> in1<3> in2<3> sl<57> vdd vss wl<3> / cell_PIM2
XI24834 bl<55> cbl<27> in1<4> in2<4> sl<55> vdd vss wl<4> / cell_PIM2
XI24183 bl<47> cbl<23> in1<25> in2<25> sl<47> vdd vss wl<25> / cell_PIM2
XI24832 bl<55> cbl<27> in1<5> in2<5> sl<55> vdd vss wl<5> / cell_PIM2
XI24831 bl<55> cbl<27> in1<6> in2<6> sl<55> vdd vss wl<6> / cell_PIM2
XI24830 bl<55> cbl<27> in1<7> in2<7> sl<55> vdd vss wl<7> / cell_PIM2
XI24833 bl<55> cbl<27> in1<3> in2<3> sl<55> vdd vss wl<3> / cell_PIM2
XI24824 bl<53> cbl<26> in1<3> in2<3> sl<53> vdd vss wl<3> / cell_PIM2
XI24173 bl<45> cbl<22> in1<26> in2<26> sl<45> vdd vss wl<26> / cell_PIM2
XI24822 bl<53> cbl<26> in1<7> in2<7> sl<53> vdd vss wl<7> / cell_PIM2
XI24821 bl<53> cbl<26> in1<6> in2<6> sl<53> vdd vss wl<6> / cell_PIM2
XI24820 bl<53> cbl<26> in1<5> in2<5> sl<53> vdd vss wl<5> / cell_PIM2
XI24823 bl<53> cbl<26> in1<4> in2<4> sl<53> vdd vss wl<4> / cell_PIM2
XI24814 bl<51> cbl<25> in1<4> in2<4> sl<51> vdd vss wl<4> / cell_PIM2
XI24163 bl<43> cbl<21> in1<25> in2<25> sl<43> vdd vss wl<25> / cell_PIM2
XI24812 bl<51> cbl<25> in1<5> in2<5> sl<51> vdd vss wl<5> / cell_PIM2
XI24811 bl<51> cbl<25> in1<6> in2<6> sl<51> vdd vss wl<6> / cell_PIM2
XI24810 bl<51> cbl<25> in1<7> in2<7> sl<51> vdd vss wl<7> / cell_PIM2
XI24813 bl<51> cbl<25> in1<3> in2<3> sl<51> vdd vss wl<3> / cell_PIM2
XI24804 bl<49> cbl<24> in1<3> in2<3> sl<49> vdd vss wl<3> / cell_PIM2
XI24153 bl<41> cbl<20> in1<25> in2<25> sl<41> vdd vss wl<25> / cell_PIM2
XI24802 bl<49> cbl<24> in1<7> in2<7> sl<49> vdd vss wl<7> / cell_PIM2
XI24801 bl<49> cbl<24> in1<6> in2<6> sl<49> vdd vss wl<6> / cell_PIM2
XI24800 bl<49> cbl<24> in1<5> in2<5> sl<49> vdd vss wl<5> / cell_PIM2
XI24803 bl<49> cbl<24> in1<4> in2<4> sl<49> vdd vss wl<4> / cell_PIM2
XI24794 bl<47> cbl<23> in1<4> in2<4> sl<47> vdd vss wl<4> / cell_PIM2
XI23018 bl<63> cbl<31> in1<61> in2<61> sl<63> vdd vss wl<61> / cell_PIM2
XI23017 bl<63> cbl<31> in1<62> in2<62> sl<63> vdd vss wl<62> / cell_PIM2
XI24222 bl<55> cbl<27> in1<26> in2<26> sl<55> vdd vss wl<26> / cell_PIM2
XI24216 bl<53> cbl<26> in1<24> in2<24> sl<53> vdd vss wl<24> / cell_PIM2
XI24215 bl<53> cbl<26> in1<23> in2<23> sl<53> vdd vss wl<23> / cell_PIM2
XI24214 bl<53> cbl<26> in1<22> in2<22> sl<53> vdd vss wl<22> / cell_PIM2
XI23568 bl<45> cbl<22> in1<43> in2<43> sl<45> vdd vss wl<43> / cell_PIM2
XI23567 bl<45> cbl<22> in1<42> in2<42> sl<45> vdd vss wl<42> / cell_PIM2
XI23566 bl<45> cbl<22> in1<41> in2<41> sl<45> vdd vss wl<41> / cell_PIM2
XI23565 bl<45> cbl<22> in1<45> in2<45> sl<45> vdd vss wl<45> / cell_PIM2
XI23564 bl<45> cbl<22> in1<44> in2<44> sl<45> vdd vss wl<44> / cell_PIM2
XI23016 bl<63> cbl<31> in1<63> in2<63> sl<63> vdd vss wl<63> / cell_PIM2
XI23015 bl<63> cbl<31> in1<64> in2<64> sl<63> vdd vss wl<64> / cell_PIM2
XI22393 bl<59> cbl<29> in1<81> in2<81> sl<59> vdd vss wl<81> / cell_PIM2
XI23010 bl<61> cbl<30> in1<62> in2<62> sl<61> vdd vss wl<62> / cell_PIM2
XI23009 bl<61> cbl<30> in1<61> in2<61> sl<61> vdd vss wl<61> / cell_PIM2
XI24212 bl<53> cbl<26> in1<25> in2<25> sl<53> vdd vss wl<25> / cell_PIM2
XI23008 bl<61> cbl<30> in1<64> in2<64> sl<61> vdd vss wl<64> / cell_PIM2
XI23007 bl<61> cbl<30> in1<63> in2<63> sl<61> vdd vss wl<63> / cell_PIM2
XI23558 bl<43> cbl<21> in1<41> in2<41> sl<43> vdd vss wl<41> / cell_PIM2
XI23557 bl<43> cbl<21> in1<42> in2<42> sl<43> vdd vss wl<42> / cell_PIM2
XI23556 bl<43> cbl<21> in1<43> in2<43> sl<43> vdd vss wl<43> / cell_PIM2
XI23555 bl<43> cbl<21> in1<44> in2<44> sl<43> vdd vss wl<44> / cell_PIM2
XI23554 bl<43> cbl<21> in1<45> in2<45> sl<43> vdd vss wl<45> / cell_PIM2
XI24206 bl<51> cbl<25> in1<22> in2<22> sl<51> vdd vss wl<22> / cell_PIM2
XI24205 bl<51> cbl<25> in1<23> in2<23> sl<51> vdd vss wl<23> / cell_PIM2
XI24204 bl<51> cbl<25> in1<24> in2<24> sl<51> vdd vss wl<24> / cell_PIM2
XI22383 bl<57> cbl<28> in1<83> in2<83> sl<57> vdd vss wl<83> / cell_PIM2
XI23002 bl<59> cbl<29> in1<61> in2<61> sl<59> vdd vss wl<61> / cell_PIM2
XI23001 bl<59> cbl<29> in1<62> in2<62> sl<59> vdd vss wl<62> / cell_PIM2
XI24202 bl<51> cbl<25> in1<26> in2<26> sl<51> vdd vss wl<26> / cell_PIM2
XI24196 bl<49> cbl<24> in1<24> in2<24> sl<49> vdd vss wl<24> / cell_PIM2
XI24195 bl<49> cbl<24> in1<23> in2<23> sl<49> vdd vss wl<23> / cell_PIM2
XI24194 bl<49> cbl<24> in1<22> in2<22> sl<49> vdd vss wl<22> / cell_PIM2
XI23548 bl<41> cbl<20> in1<41> in2<41> sl<41> vdd vss wl<41> / cell_PIM2
XI23547 bl<41> cbl<20> in1<42> in2<42> sl<41> vdd vss wl<42> / cell_PIM2
XI23546 bl<41> cbl<20> in1<43> in2<43> sl<41> vdd vss wl<43> / cell_PIM2
XI23545 bl<41> cbl<20> in1<44> in2<44> sl<41> vdd vss wl<44> / cell_PIM2
XI23544 bl<41> cbl<20> in1<45> in2<45> sl<41> vdd vss wl<45> / cell_PIM2
XI23000 bl<59> cbl<29> in1<63> in2<63> sl<59> vdd vss wl<63> / cell_PIM2
XI22999 bl<59> cbl<29> in1<64> in2<64> sl<59> vdd vss wl<64> / cell_PIM2
XI22378 bl<55> cbl<27> in1<80> in2<80> sl<55> vdd vss wl<80> / cell_PIM2
XI22994 bl<57> cbl<28> in1<61> in2<61> sl<57> vdd vss wl<61> / cell_PIM2
XI22993 bl<57> cbl<28> in1<62> in2<62> sl<57> vdd vss wl<62> / cell_PIM2
XI24192 bl<49> cbl<24> in1<25> in2<25> sl<49> vdd vss wl<25> / cell_PIM2
XI22368 bl<53> cbl<26> in1<83> in2<83> sl<53> vdd vss wl<83> / cell_PIM2
XI22992 bl<57> cbl<28> in1<63> in2<63> sl<57> vdd vss wl<63> / cell_PIM2
XI22991 bl<57> cbl<28> in1<64> in2<64> sl<57> vdd vss wl<64> / cell_PIM2
XI23538 bl<39> cbl<19> in1<41> in2<41> sl<39> vdd vss wl<41> / cell_PIM2
XI23537 bl<39> cbl<19> in1<42> in2<42> sl<39> vdd vss wl<42> / cell_PIM2
XI23536 bl<39> cbl<19> in1<43> in2<43> sl<39> vdd vss wl<43> / cell_PIM2
XI23535 bl<39> cbl<19> in1<44> in2<44> sl<39> vdd vss wl<44> / cell_PIM2
XI23534 bl<39> cbl<19> in1<45> in2<45> sl<39> vdd vss wl<45> / cell_PIM2
XI24186 bl<47> cbl<23> in1<22> in2<22> sl<47> vdd vss wl<22> / cell_PIM2
XI24185 bl<47> cbl<23> in1<23> in2<23> sl<47> vdd vss wl<23> / cell_PIM2
XI24184 bl<47> cbl<23> in1<24> in2<24> sl<47> vdd vss wl<24> / cell_PIM2
XI22986 bl<55> cbl<27> in1<61> in2<61> sl<55> vdd vss wl<61> / cell_PIM2
XI22985 bl<55> cbl<27> in1<62> in2<62> sl<55> vdd vss wl<62> / cell_PIM2
XI24182 bl<47> cbl<23> in1<26> in2<26> sl<47> vdd vss wl<26> / cell_PIM2
XI24176 bl<45> cbl<22> in1<24> in2<24> sl<45> vdd vss wl<24> / cell_PIM2
XI24175 bl<45> cbl<22> in1<23> in2<23> sl<45> vdd vss wl<23> / cell_PIM2
XI24174 bl<45> cbl<22> in1<22> in2<22> sl<45> vdd vss wl<22> / cell_PIM2
XI23528 bl<37> cbl<18> in1<43> in2<43> sl<37> vdd vss wl<43> / cell_PIM2
XI23527 bl<37> cbl<18> in1<42> in2<42> sl<37> vdd vss wl<42> / cell_PIM2
XI23526 bl<37> cbl<18> in1<41> in2<41> sl<37> vdd vss wl<41> / cell_PIM2
XI23525 bl<37> cbl<18> in1<45> in2<45> sl<37> vdd vss wl<45> / cell_PIM2
XI23524 bl<37> cbl<18> in1<44> in2<44> sl<37> vdd vss wl<44> / cell_PIM2
XI22984 bl<55> cbl<27> in1<63> in2<63> sl<55> vdd vss wl<63> / cell_PIM2
XI22983 bl<55> cbl<27> in1<64> in2<64> sl<55> vdd vss wl<64> / cell_PIM2
XI22353 bl<49> cbl<24> in1<80> in2<80> sl<49> vdd vss wl<80> / cell_PIM2
XI22978 bl<53> cbl<26> in1<62> in2<62> sl<53> vdd vss wl<62> / cell_PIM2
XI22977 bl<53> cbl<26> in1<61> in2<61> sl<53> vdd vss wl<61> / cell_PIM2
XI24172 bl<45> cbl<22> in1<25> in2<25> sl<45> vdd vss wl<25> / cell_PIM2
XI22976 bl<53> cbl<26> in1<64> in2<64> sl<53> vdd vss wl<64> / cell_PIM2
XI22975 bl<53> cbl<26> in1<63> in2<63> sl<53> vdd vss wl<63> / cell_PIM2
XI23518 bl<35> cbl<17> in1<41> in2<41> sl<35> vdd vss wl<41> / cell_PIM2
XI23517 bl<35> cbl<17> in1<42> in2<42> sl<35> vdd vss wl<42> / cell_PIM2
XI23516 bl<35> cbl<17> in1<43> in2<43> sl<35> vdd vss wl<43> / cell_PIM2
XI23515 bl<35> cbl<17> in1<44> in2<44> sl<35> vdd vss wl<44> / cell_PIM2
XI23514 bl<35> cbl<17> in1<45> in2<45> sl<35> vdd vss wl<45> / cell_PIM2
XI24166 bl<43> cbl<21> in1<22> in2<22> sl<43> vdd vss wl<22> / cell_PIM2
XI24165 bl<43> cbl<21> in1<23> in2<23> sl<43> vdd vss wl<23> / cell_PIM2
XI24164 bl<43> cbl<21> in1<24> in2<24> sl<43> vdd vss wl<24> / cell_PIM2
XI22343 bl<47> cbl<23> in1<83> in2<83> sl<47> vdd vss wl<83> / cell_PIM2
XI22970 bl<51> cbl<25> in1<61> in2<61> sl<51> vdd vss wl<61> / cell_PIM2
XI22969 bl<51> cbl<25> in1<62> in2<62> sl<51> vdd vss wl<62> / cell_PIM2
XI24162 bl<43> cbl<21> in1<26> in2<26> sl<43> vdd vss wl<26> / cell_PIM2
XI24156 bl<41> cbl<20> in1<22> in2<22> sl<41> vdd vss wl<22> / cell_PIM2
XI24155 bl<41> cbl<20> in1<23> in2<23> sl<41> vdd vss wl<23> / cell_PIM2
XI24154 bl<41> cbl<20> in1<24> in2<24> sl<41> vdd vss wl<24> / cell_PIM2
XI23508 bl<33> cbl<16> in1<43> in2<43> sl<33> vdd vss wl<43> / cell_PIM2
XI23507 bl<33> cbl<16> in1<42> in2<42> sl<33> vdd vss wl<42> / cell_PIM2
XI23506 bl<33> cbl<16> in1<41> in2<41> sl<33> vdd vss wl<41> / cell_PIM2
XI23505 bl<33> cbl<16> in1<45> in2<45> sl<33> vdd vss wl<45> / cell_PIM2
XI23504 bl<33> cbl<16> in1<44> in2<44> sl<33> vdd vss wl<44> / cell_PIM2
XI22968 bl<51> cbl<25> in1<63> in2<63> sl<51> vdd vss wl<63> / cell_PIM2
XI22967 bl<51> cbl<25> in1<64> in2<64> sl<51> vdd vss wl<64> / cell_PIM2
XI22338 bl<45> cbl<22> in1<81> in2<81> sl<45> vdd vss wl<81> / cell_PIM2
XI22962 bl<49> cbl<24> in1<62> in2<62> sl<49> vdd vss wl<62> / cell_PIM2
XI22961 bl<49> cbl<24> in1<61> in2<61> sl<49> vdd vss wl<61> / cell_PIM2
XI24152 bl<41> cbl<20> in1<26> in2<26> sl<41> vdd vss wl<26> / cell_PIM2
XI22328 bl<43> cbl<21> in1<82> in2<82> sl<43> vdd vss wl<82> / cell_PIM2
XI22960 bl<49> cbl<24> in1<64> in2<64> sl<49> vdd vss wl<64> / cell_PIM2
XI22959 bl<49> cbl<24> in1<63> in2<63> sl<49> vdd vss wl<63> / cell_PIM2
XI23498 bl<63> cbl<31> in1<46> in2<46> sl<63> vdd vss wl<46> / cell_PIM2
XI23497 bl<63> cbl<31> in1<47> in2<47> sl<63> vdd vss wl<47> / cell_PIM2
XI23496 bl<63> cbl<31> in1<48> in2<48> sl<63> vdd vss wl<48> / cell_PIM2
XI23495 bl<63> cbl<31> in1<49> in2<49> sl<63> vdd vss wl<49> / cell_PIM2
XI23494 bl<63> cbl<31> in1<50> in2<50> sl<63> vdd vss wl<50> / cell_PIM2
XI24146 bl<39> cbl<19> in1<22> in2<22> sl<39> vdd vss wl<22> / cell_PIM2
XI24145 bl<39> cbl<19> in1<23> in2<23> sl<39> vdd vss wl<23> / cell_PIM2
XI24144 bl<39> cbl<19> in1<24> in2<24> sl<39> vdd vss wl<24> / cell_PIM2
XI21103 bl<45> cbl<22> in1<118> in2<118> sl<45> vdd vss wl<118> / cell_PIM2
XI21102 bl<45> cbl<22> in1<122> in2<122> sl<45> vdd vss wl<122> / cell_PIM2
XI21101 bl<45> cbl<22> in1<121> in2<121> sl<45> vdd vss wl<121> / cell_PIM2
XI21100 bl<45> cbl<22> in1<120> in2<120> sl<45> vdd vss wl<120> / cell_PIM2
XI21752 bl<53> cbl<26> in1<100> in2<100> sl<53> vdd vss wl<100> / cell_PIM2
XI21751 bl<53> cbl<26> in1<99> in2<99> sl<53> vdd vss wl<99> / cell_PIM2
XI21750 bl<53> cbl<26> in1<103> in2<103> sl<53> vdd vss wl<103> / cell_PIM2
XI21749 bl<53> cbl<26> in1<102> in2<102> sl<53> vdd vss wl<102> / cell_PIM2
XI22402 bl<61> cbl<30> in1<81> in2<81> sl<61> vdd vss wl<81> / cell_PIM2
XI22401 bl<61> cbl<30> in1<80> in2<80> sl<61> vdd vss wl<80> / cell_PIM2
XI22400 bl<61> cbl<30> in1<83> in2<83> sl<61> vdd vss wl<83> / cell_PIM2
XI22399 bl<61> cbl<30> in1<82> in2<82> sl<61> vdd vss wl<82> / cell_PIM2
XI21748 bl<53> cbl<26> in1<101> in2<101> sl<53> vdd vss wl<101> / cell_PIM2
XI21094 bl<43> cbl<21> in1<118> in2<118> sl<43> vdd vss wl<118> / cell_PIM2
XI22394 bl<59> cbl<29> in1<80> in2<80> sl<59> vdd vss wl<80> / cell_PIM2
XI21093 bl<43> cbl<21> in1<119> in2<119> sl<43> vdd vss wl<119> / cell_PIM2
XI21092 bl<43> cbl<21> in1<120> in2<120> sl<43> vdd vss wl<120> / cell_PIM2
XI21091 bl<43> cbl<21> in1<121> in2<121> sl<43> vdd vss wl<121> / cell_PIM2
XI21090 bl<43> cbl<21> in1<122> in2<122> sl<43> vdd vss wl<122> / cell_PIM2
XI21742 bl<51> cbl<25> in1<99> in2<99> sl<51> vdd vss wl<99> / cell_PIM2
XI21741 bl<51> cbl<25> in1<100> in2<100> sl<51> vdd vss wl<100> / cell_PIM2
XI21740 bl<51> cbl<25> in1<101> in2<101> sl<51> vdd vss wl<101> / cell_PIM2
XI21739 bl<51> cbl<25> in1<102> in2<102> sl<51> vdd vss wl<102> / cell_PIM2
XI22392 bl<59> cbl<29> in1<82> in2<82> sl<59> vdd vss wl<82> / cell_PIM2
XI22391 bl<59> cbl<29> in1<83> in2<83> sl<59> vdd vss wl<83> / cell_PIM2
XI21084 bl<41> cbl<20> in1<118> in2<118> sl<41> vdd vss wl<118> / cell_PIM2
XI21738 bl<51> cbl<25> in1<103> in2<103> sl<51> vdd vss wl<103> / cell_PIM2
XI22386 bl<57> cbl<28> in1<80> in2<80> sl<57> vdd vss wl<80> / cell_PIM2
XI22385 bl<57> cbl<28> in1<81> in2<81> sl<57> vdd vss wl<81> / cell_PIM2
XI22384 bl<57> cbl<28> in1<82> in2<82> sl<57> vdd vss wl<82> / cell_PIM2
XI21083 bl<41> cbl<20> in1<119> in2<119> sl<41> vdd vss wl<119> / cell_PIM2
XI21082 bl<41> cbl<20> in1<120> in2<120> sl<41> vdd vss wl<120> / cell_PIM2
XI21081 bl<41> cbl<20> in1<121> in2<121> sl<41> vdd vss wl<121> / cell_PIM2
XI21080 bl<41> cbl<20> in1<122> in2<122> sl<41> vdd vss wl<122> / cell_PIM2
XI21732 bl<49> cbl<24> in1<100> in2<100> sl<49> vdd vss wl<100> / cell_PIM2
XI21731 bl<49> cbl<24> in1<99> in2<99> sl<49> vdd vss wl<99> / cell_PIM2
XI21730 bl<49> cbl<24> in1<103> in2<103> sl<49> vdd vss wl<103> / cell_PIM2
XI21729 bl<49> cbl<24> in1<102> in2<102> sl<49> vdd vss wl<102> / cell_PIM2
XI22377 bl<55> cbl<27> in1<81> in2<81> sl<55> vdd vss wl<81> / cell_PIM2
XI22376 bl<55> cbl<27> in1<82> in2<82> sl<55> vdd vss wl<82> / cell_PIM2
XI22375 bl<55> cbl<27> in1<83> in2<83> sl<55> vdd vss wl<83> / cell_PIM2
XI21728 bl<49> cbl<24> in1<101> in2<101> sl<49> vdd vss wl<101> / cell_PIM2
XI21074 bl<39> cbl<19> in1<118> in2<118> sl<39> vdd vss wl<118> / cell_PIM2
XI21073 bl<39> cbl<19> in1<119> in2<119> sl<39> vdd vss wl<119> / cell_PIM2
XI21072 bl<39> cbl<19> in1<120> in2<120> sl<39> vdd vss wl<120> / cell_PIM2
XI21071 bl<39> cbl<19> in1<121> in2<121> sl<39> vdd vss wl<121> / cell_PIM2
XI21070 bl<39> cbl<19> in1<122> in2<122> sl<39> vdd vss wl<122> / cell_PIM2
XI21722 bl<47> cbl<23> in1<99> in2<99> sl<47> vdd vss wl<99> / cell_PIM2
XI21721 bl<47> cbl<23> in1<100> in2<100> sl<47> vdd vss wl<100> / cell_PIM2
XI21720 bl<47> cbl<23> in1<101> in2<101> sl<47> vdd vss wl<101> / cell_PIM2
XI21719 bl<47> cbl<23> in1<102> in2<102> sl<47> vdd vss wl<102> / cell_PIM2
XI22370 bl<53> cbl<26> in1<81> in2<81> sl<53> vdd vss wl<81> / cell_PIM2
XI22369 bl<53> cbl<26> in1<80> in2<80> sl<53> vdd vss wl<80> / cell_PIM2
XI21064 bl<37> cbl<18> in1<119> in2<119> sl<37> vdd vss wl<119> / cell_PIM2
XI21718 bl<47> cbl<23> in1<103> in2<103> sl<47> vdd vss wl<103> / cell_PIM2
XI22367 bl<53> cbl<26> in1<82> in2<82> sl<53> vdd vss wl<82> / cell_PIM2
XI21063 bl<37> cbl<18> in1<118> in2<118> sl<37> vdd vss wl<118> / cell_PIM2
XI21062 bl<37> cbl<18> in1<122> in2<122> sl<37> vdd vss wl<122> / cell_PIM2
XI21061 bl<37> cbl<18> in1<121> in2<121> sl<37> vdd vss wl<121> / cell_PIM2
XI21060 bl<37> cbl<18> in1<120> in2<120> sl<37> vdd vss wl<120> / cell_PIM2
XI21712 bl<45> cbl<22> in1<100> in2<100> sl<45> vdd vss wl<100> / cell_PIM2
XI21711 bl<45> cbl<22> in1<99> in2<99> sl<45> vdd vss wl<99> / cell_PIM2
XI21710 bl<45> cbl<22> in1<103> in2<103> sl<45> vdd vss wl<103> / cell_PIM2
XI21709 bl<45> cbl<22> in1<102> in2<102> sl<45> vdd vss wl<102> / cell_PIM2
XI22362 bl<51> cbl<25> in1<80> in2<80> sl<51> vdd vss wl<80> / cell_PIM2
XI22361 bl<51> cbl<25> in1<81> in2<81> sl<51> vdd vss wl<81> / cell_PIM2
XI22360 bl<51> cbl<25> in1<82> in2<82> sl<51> vdd vss wl<82> / cell_PIM2
XI22359 bl<51> cbl<25> in1<83> in2<83> sl<51> vdd vss wl<83> / cell_PIM2
XI21708 bl<45> cbl<22> in1<101> in2<101> sl<45> vdd vss wl<101> / cell_PIM2
XI21054 bl<35> cbl<17> in1<118> in2<118> sl<35> vdd vss wl<118> / cell_PIM2
XI22354 bl<49> cbl<24> in1<81> in2<81> sl<49> vdd vss wl<81> / cell_PIM2
XI21053 bl<35> cbl<17> in1<119> in2<119> sl<35> vdd vss wl<119> / cell_PIM2
XI21052 bl<35> cbl<17> in1<120> in2<120> sl<35> vdd vss wl<120> / cell_PIM2
XI21051 bl<35> cbl<17> in1<121> in2<121> sl<35> vdd vss wl<121> / cell_PIM2
XI21050 bl<35> cbl<17> in1<122> in2<122> sl<35> vdd vss wl<122> / cell_PIM2
XI21702 bl<43> cbl<21> in1<99> in2<99> sl<43> vdd vss wl<99> / cell_PIM2
XI21701 bl<43> cbl<21> in1<100> in2<100> sl<43> vdd vss wl<100> / cell_PIM2
XI21700 bl<43> cbl<21> in1<101> in2<101> sl<43> vdd vss wl<101> / cell_PIM2
XI21699 bl<43> cbl<21> in1<102> in2<102> sl<43> vdd vss wl<102> / cell_PIM2
XI22352 bl<49> cbl<24> in1<83> in2<83> sl<49> vdd vss wl<83> / cell_PIM2
XI22351 bl<49> cbl<24> in1<82> in2<82> sl<49> vdd vss wl<82> / cell_PIM2
XI21044 bl<33> cbl<16> in1<119> in2<119> sl<33> vdd vss wl<119> / cell_PIM2
XI21698 bl<43> cbl<21> in1<103> in2<103> sl<43> vdd vss wl<103> / cell_PIM2
XI22346 bl<47> cbl<23> in1<80> in2<80> sl<47> vdd vss wl<80> / cell_PIM2
XI22345 bl<47> cbl<23> in1<81> in2<81> sl<47> vdd vss wl<81> / cell_PIM2
XI22344 bl<47> cbl<23> in1<82> in2<82> sl<47> vdd vss wl<82> / cell_PIM2
XI21043 bl<33> cbl<16> in1<118> in2<118> sl<33> vdd vss wl<118> / cell_PIM2
XI21042 bl<33> cbl<16> in1<122> in2<122> sl<33> vdd vss wl<122> / cell_PIM2
XI21041 bl<33> cbl<16> in1<121> in2<121> sl<33> vdd vss wl<121> / cell_PIM2
XI21040 bl<33> cbl<16> in1<120> in2<120> sl<33> vdd vss wl<120> / cell_PIM2
XI21692 bl<41> cbl<20> in1<99> in2<99> sl<41> vdd vss wl<99> / cell_PIM2
XI21691 bl<41> cbl<20> in1<100> in2<100> sl<41> vdd vss wl<100> / cell_PIM2
XI21690 bl<41> cbl<20> in1<101> in2<101> sl<41> vdd vss wl<101> / cell_PIM2
XI21689 bl<41> cbl<20> in1<102> in2<102> sl<41> vdd vss wl<102> / cell_PIM2
XI22337 bl<45> cbl<22> in1<80> in2<80> sl<45> vdd vss wl<80> / cell_PIM2
XI22336 bl<45> cbl<22> in1<83> in2<83> sl<45> vdd vss wl<83> / cell_PIM2
XI22335 bl<45> cbl<22> in1<82> in2<82> sl<45> vdd vss wl<82> / cell_PIM2
XI21688 bl<41> cbl<20> in1<103> in2<103> sl<41> vdd vss wl<103> / cell_PIM2
XI21034 bl<63> cbl<31> in1<127> in2<127> sl<63> vdd vss wl<127> / cell_PIM2
XI21033 bl<63> cbl<31> in1<126> in2<126> sl<63> vdd vss wl<126> / cell_PIM2
XI21032 bl<63> cbl<31> in1<125> in2<125> sl<63> vdd vss wl<125> / cell_PIM2
XI21031 bl<63> cbl<31> in1<123> in2<123> sl<63> vdd vss wl<123> / cell_PIM2
XI21030 bl<63> cbl<31> in1<124> in2<124> sl<63> vdd vss wl<124> / cell_PIM2
XI21682 bl<39> cbl<19> in1<99> in2<99> sl<39> vdd vss wl<99> / cell_PIM2
XI21681 bl<39> cbl<19> in1<100> in2<100> sl<39> vdd vss wl<100> / cell_PIM2
XI21680 bl<39> cbl<19> in1<101> in2<101> sl<39> vdd vss wl<101> / cell_PIM2
XI21679 bl<39> cbl<19> in1<102> in2<102> sl<39> vdd vss wl<102> / cell_PIM2
XI22330 bl<43> cbl<21> in1<80> in2<80> sl<43> vdd vss wl<80> / cell_PIM2
XI22329 bl<43> cbl<21> in1<81> in2<81> sl<43> vdd vss wl<81> / cell_PIM2
XI21024 bl<61> cbl<30> in1<127> in2<127> sl<61> vdd vss wl<127> / cell_PIM2
XI21678 bl<39> cbl<19> in1<103> in2<103> sl<39> vdd vss wl<103> / cell_PIM2
XI22327 bl<43> cbl<21> in1<83> in2<83> sl<43> vdd vss wl<83> / cell_PIM2
XI19280 bl<29> cbl<14> in1<100> in2<100> sl<29> vdd vss wl<100> / cell_PIM2
XI19279 bl<29> cbl<14> in1<99> in2<99> sl<29> vdd vss wl<99> / cell_PIM2
XI19898 bl<31> cbl<15> in1<61> in2<61> sl<31> vdd vss wl<61> / cell_PIM2
XI19897 bl<31> cbl<15> in1<62> in2<62> sl<31> vdd vss wl<62> / cell_PIM2
XI20452 bl<17> cbl<8> in1<24> in2<24> sl<17> vdd vss wl<24> / cell_PIM2
XI20451 bl<17> cbl<8> in1<23> in2<23> sl<17> vdd vss wl<23> / cell_PIM2
XI20450 bl<17> cbl<8> in1<22> in2<22> sl<17> vdd vss wl<22> / cell_PIM2
XI20449 bl<17> cbl<8> in1<26> in2<26> sl<17> vdd vss wl<26> / cell_PIM2
XI20448 bl<17> cbl<8> in1<25> in2<25> sl<17> vdd vss wl<25> / cell_PIM2
XI19896 bl<31> cbl<15> in1<63> in2<63> sl<31> vdd vss wl<63> / cell_PIM2
XI19895 bl<31> cbl<15> in1<64> in2<64> sl<31> vdd vss wl<64> / cell_PIM2
XI19278 bl<29> cbl<14> in1<103> in2<103> sl<29> vdd vss wl<103> / cell_PIM2
XI19277 bl<29> cbl<14> in1<102> in2<102> sl<29> vdd vss wl<102> / cell_PIM2
XI19276 bl<29> cbl<14> in1<101> in2<101> sl<29> vdd vss wl<101> / cell_PIM2
XI19270 bl<27> cbl<13> in1<99> in2<99> sl<27> vdd vss wl<99> / cell_PIM2
XI19269 bl<27> cbl<13> in1<100> in2<100> sl<27> vdd vss wl<100> / cell_PIM2
XI19890 bl<29> cbl<14> in1<62> in2<62> sl<29> vdd vss wl<62> / cell_PIM2
XI19889 bl<29> cbl<14> in1<61> in2<61> sl<29> vdd vss wl<61> / cell_PIM2
XI20442 bl<31> cbl<15> in1<27> in2<27> sl<31> vdd vss wl<27> / cell_PIM2
XI20441 bl<31> cbl<15> in1<28> in2<28> sl<31> vdd vss wl<28> / cell_PIM2
XI20440 bl<31> cbl<15> in1<29> in2<29> sl<31> vdd vss wl<29> / cell_PIM2
XI20439 bl<31> cbl<15> in1<30> in2<30> sl<31> vdd vss wl<30> / cell_PIM2
XI19267 bl<27> cbl<13> in1<102> in2<102> sl<27> vdd vss wl<102> / cell_PIM2
XI19266 bl<27> cbl<13> in1<103> in2<103> sl<27> vdd vss wl<103> / cell_PIM2
XI19268 bl<27> cbl<13> in1<101> in2<101> sl<27> vdd vss wl<101> / cell_PIM2
XI19888 bl<29> cbl<14> in1<64> in2<64> sl<29> vdd vss wl<64> / cell_PIM2
XI19887 bl<29> cbl<14> in1<63> in2<63> sl<29> vdd vss wl<63> / cell_PIM2
XI20438 bl<31> cbl<15> in1<31> in2<31> sl<31> vdd vss wl<31> / cell_PIM2
XI19260 bl<25> cbl<12> in1<99> in2<99> sl<25> vdd vss wl<99> / cell_PIM2
XI19259 bl<25> cbl<12> in1<100> in2<100> sl<25> vdd vss wl<100> / cell_PIM2
XI19882 bl<27> cbl<13> in1<61> in2<61> sl<27> vdd vss wl<61> / cell_PIM2
XI19881 bl<27> cbl<13> in1<62> in2<62> sl<27> vdd vss wl<62> / cell_PIM2
XI20432 bl<29> cbl<14> in1<28> in2<28> sl<29> vdd vss wl<28> / cell_PIM2
XI20431 bl<29> cbl<14> in1<27> in2<27> sl<29> vdd vss wl<27> / cell_PIM2
XI20430 bl<29> cbl<14> in1<31> in2<31> sl<29> vdd vss wl<31> / cell_PIM2
XI20429 bl<29> cbl<14> in1<30> in2<30> sl<29> vdd vss wl<30> / cell_PIM2
XI20428 bl<29> cbl<14> in1<29> in2<29> sl<29> vdd vss wl<29> / cell_PIM2
XI19880 bl<27> cbl<13> in1<63> in2<63> sl<27> vdd vss wl<63> / cell_PIM2
XI19879 bl<27> cbl<13> in1<64> in2<64> sl<27> vdd vss wl<64> / cell_PIM2
XI19258 bl<25> cbl<12> in1<101> in2<101> sl<25> vdd vss wl<101> / cell_PIM2
XI19257 bl<25> cbl<12> in1<102> in2<102> sl<25> vdd vss wl<102> / cell_PIM2
XI19256 bl<25> cbl<12> in1<103> in2<103> sl<25> vdd vss wl<103> / cell_PIM2
XI19250 bl<23> cbl<11> in1<99> in2<99> sl<23> vdd vss wl<99> / cell_PIM2
XI19249 bl<23> cbl<11> in1<100> in2<100> sl<23> vdd vss wl<100> / cell_PIM2
XI19874 bl<25> cbl<12> in1<61> in2<61> sl<25> vdd vss wl<61> / cell_PIM2
XI19873 bl<25> cbl<12> in1<62> in2<62> sl<25> vdd vss wl<62> / cell_PIM2
XI20422 bl<27> cbl<13> in1<27> in2<27> sl<27> vdd vss wl<27> / cell_PIM2
XI20421 bl<27> cbl<13> in1<28> in2<28> sl<27> vdd vss wl<28> / cell_PIM2
XI20420 bl<27> cbl<13> in1<29> in2<29> sl<27> vdd vss wl<29> / cell_PIM2
XI20419 bl<27> cbl<13> in1<30> in2<30> sl<27> vdd vss wl<30> / cell_PIM2
XI19247 bl<23> cbl<11> in1<102> in2<102> sl<23> vdd vss wl<102> / cell_PIM2
XI19246 bl<23> cbl<11> in1<103> in2<103> sl<23> vdd vss wl<103> / cell_PIM2
XI19248 bl<23> cbl<11> in1<101> in2<101> sl<23> vdd vss wl<101> / cell_PIM2
XI19872 bl<25> cbl<12> in1<63> in2<63> sl<25> vdd vss wl<63> / cell_PIM2
XI19871 bl<25> cbl<12> in1<64> in2<64> sl<25> vdd vss wl<64> / cell_PIM2
XI20418 bl<27> cbl<13> in1<31> in2<31> sl<27> vdd vss wl<31> / cell_PIM2
XI19240 bl<21> cbl<10> in1<100> in2<100> sl<21> vdd vss wl<100> / cell_PIM2
XI19239 bl<21> cbl<10> in1<99> in2<99> sl<21> vdd vss wl<99> / cell_PIM2
XI19866 bl<23> cbl<11> in1<61> in2<61> sl<23> vdd vss wl<61> / cell_PIM2
XI19865 bl<23> cbl<11> in1<62> in2<62> sl<23> vdd vss wl<62> / cell_PIM2
XI20412 bl<25> cbl<12> in1<27> in2<27> sl<25> vdd vss wl<27> / cell_PIM2
XI20411 bl<25> cbl<12> in1<28> in2<28> sl<25> vdd vss wl<28> / cell_PIM2
XI20410 bl<25> cbl<12> in1<29> in2<29> sl<25> vdd vss wl<29> / cell_PIM2
XI20409 bl<25> cbl<12> in1<30> in2<30> sl<25> vdd vss wl<30> / cell_PIM2
XI20408 bl<25> cbl<12> in1<31> in2<31> sl<25> vdd vss wl<31> / cell_PIM2
XI19864 bl<23> cbl<11> in1<63> in2<63> sl<23> vdd vss wl<63> / cell_PIM2
XI19863 bl<23> cbl<11> in1<64> in2<64> sl<23> vdd vss wl<64> / cell_PIM2
XI19238 bl<21> cbl<10> in1<103> in2<103> sl<21> vdd vss wl<103> / cell_PIM2
XI19237 bl<21> cbl<10> in1<102> in2<102> sl<21> vdd vss wl<102> / cell_PIM2
XI19236 bl<21> cbl<10> in1<101> in2<101> sl<21> vdd vss wl<101> / cell_PIM2
XI19230 bl<19> cbl<9> in1<99> in2<99> sl<19> vdd vss wl<99> / cell_PIM2
XI19229 bl<19> cbl<9> in1<100> in2<100> sl<19> vdd vss wl<100> / cell_PIM2
XI19858 bl<21> cbl<10> in1<62> in2<62> sl<21> vdd vss wl<62> / cell_PIM2
XI19857 bl<21> cbl<10> in1<61> in2<61> sl<21> vdd vss wl<61> / cell_PIM2
XI20402 bl<23> cbl<11> in1<27> in2<27> sl<23> vdd vss wl<27> / cell_PIM2
XI20401 bl<23> cbl<11> in1<28> in2<28> sl<23> vdd vss wl<28> / cell_PIM2
XI20400 bl<23> cbl<11> in1<29> in2<29> sl<23> vdd vss wl<29> / cell_PIM2
XI20399 bl<23> cbl<11> in1<30> in2<30> sl<23> vdd vss wl<30> / cell_PIM2
XI19227 bl<19> cbl<9> in1<102> in2<102> sl<19> vdd vss wl<102> / cell_PIM2
XI19226 bl<19> cbl<9> in1<103> in2<103> sl<19> vdd vss wl<103> / cell_PIM2
XI19228 bl<19> cbl<9> in1<101> in2<101> sl<19> vdd vss wl<101> / cell_PIM2
XI19856 bl<21> cbl<10> in1<64> in2<64> sl<21> vdd vss wl<64> / cell_PIM2
XI19855 bl<21> cbl<10> in1<63> in2<63> sl<21> vdd vss wl<63> / cell_PIM2
XI20398 bl<23> cbl<11> in1<31> in2<31> sl<23> vdd vss wl<31> / cell_PIM2
XI19220 bl<17> cbl<8> in1<100> in2<100> sl<17> vdd vss wl<100> / cell_PIM2
XI19219 bl<17> cbl<8> in1<99> in2<99> sl<17> vdd vss wl<99> / cell_PIM2
XI19850 bl<19> cbl<9> in1<61> in2<61> sl<19> vdd vss wl<61> / cell_PIM2
XI19849 bl<19> cbl<9> in1<62> in2<62> sl<19> vdd vss wl<62> / cell_PIM2
XI20392 bl<21> cbl<10> in1<28> in2<28> sl<21> vdd vss wl<28> / cell_PIM2
XI20391 bl<21> cbl<10> in1<27> in2<27> sl<21> vdd vss wl<27> / cell_PIM2
XI20390 bl<21> cbl<10> in1<31> in2<31> sl<21> vdd vss wl<31> / cell_PIM2
XI20389 bl<21> cbl<10> in1<30> in2<30> sl<21> vdd vss wl<30> / cell_PIM2
XI20388 bl<21> cbl<10> in1<29> in2<29> sl<21> vdd vss wl<29> / cell_PIM2
XI19848 bl<19> cbl<9> in1<63> in2<63> sl<19> vdd vss wl<63> / cell_PIM2
XI19847 bl<19> cbl<9> in1<64> in2<64> sl<19> vdd vss wl<64> / cell_PIM2
XI19218 bl<17> cbl<8> in1<103> in2<103> sl<17> vdd vss wl<103> / cell_PIM2
XI19217 bl<17> cbl<8> in1<102> in2<102> sl<17> vdd vss wl<102> / cell_PIM2
XI19216 bl<17> cbl<8> in1<101> in2<101> sl<17> vdd vss wl<101> / cell_PIM2
XI19210 bl<31> cbl<15> in1<104> in2<104> sl<31> vdd vss wl<104> / cell_PIM2
XI19209 bl<31> cbl<15> in1<105> in2<105> sl<31> vdd vss wl<105> / cell_PIM2
XI19842 bl<17> cbl<8> in1<62> in2<62> sl<17> vdd vss wl<62> / cell_PIM2
XI19841 bl<17> cbl<8> in1<61> in2<61> sl<17> vdd vss wl<61> / cell_PIM2
XI20382 bl<19> cbl<9> in1<27> in2<27> sl<19> vdd vss wl<27> / cell_PIM2
XI20381 bl<19> cbl<9> in1<28> in2<28> sl<19> vdd vss wl<28> / cell_PIM2
XI20380 bl<19> cbl<9> in1<29> in2<29> sl<19> vdd vss wl<29> / cell_PIM2
XI20379 bl<19> cbl<9> in1<30> in2<30> sl<19> vdd vss wl<30> / cell_PIM2
XI19207 bl<31> cbl<15> in1<107> in2<107> sl<31> vdd vss wl<107> / cell_PIM2
XI19208 bl<31> cbl<15> in1<106> in2<106> sl<31> vdd vss wl<106> / cell_PIM2
XI19840 bl<17> cbl<8> in1<64> in2<64> sl<17> vdd vss wl<64> / cell_PIM2
XI19839 bl<17> cbl<8> in1<63> in2<63> sl<17> vdd vss wl<63> / cell_PIM2
XI20378 bl<19> cbl<9> in1<31> in2<31> sl<19> vdd vss wl<31> / cell_PIM2
XI17330 bl<5> cbl<2> in1<119> in2<119> sl<5> vdd vss wl<119> / cell_PIM2
XI17329 bl<5> cbl<2> in1<118> in2<118> sl<5> vdd vss wl<118> / cell_PIM2
XI18633 bl<9> cbl<4> in1<21> in2<21> sl<9> vdd vss wl<21> / cell_PIM2
XI18632 bl<9> cbl<4> in1<20> in2<20> sl<9> vdd vss wl<20> / cell_PIM2
XI18626 bl<15> cbl<7> in1<25> in2<25> sl<15> vdd vss wl<25> / cell_PIM2
XI18625 bl<15> cbl<7> in1<26> in2<26> sl<15> vdd vss wl<26> / cell_PIM2
XI18624 bl<15> cbl<7> in1<27> in2<27> sl<15> vdd vss wl<27> / cell_PIM2
XI17978 bl<15> cbl<7> in1<106> in2<106> sl<15> vdd vss wl<106> / cell_PIM2
XI17977 bl<15> cbl<7> in1<107> in2<107> sl<15> vdd vss wl<107> / cell_PIM2
XI17976 bl<15> cbl<7> in1<108> in2<108> sl<15> vdd vss wl<108> / cell_PIM2
XI17975 bl<15> cbl<7> in1<109> in2<109> sl<15> vdd vss wl<109> / cell_PIM2
XI17974 bl<15> cbl<7> in1<110> in2<110> sl<15> vdd vss wl<110> / cell_PIM2
XI17328 bl<5> cbl<2> in1<117> in2<117> sl<5> vdd vss wl<117> / cell_PIM2
XI17327 bl<5> cbl<2> in1<116> in2<116> sl<5> vdd vss wl<116> / cell_PIM2
XI17322 bl<7> cbl<3> in1<120> in2<120> sl<7> vdd vss wl<120> / cell_PIM2
XI17321 bl<7> cbl<3> in1<121> in2<121> sl<7> vdd vss wl<121> / cell_PIM2
XI17320 bl<7> cbl<3> in1<122> in2<122> sl<7> vdd vss wl<122> / cell_PIM2
XI17319 bl<7> cbl<3> in1<123> in2<123> sl<7> vdd vss wl<123> / cell_PIM2
XI18623 bl<15> cbl<7> in1<28> in2<28> sl<15> vdd vss wl<28> / cell_PIM2
XI17318 bl<7> cbl<3> in1<124> in2<124> sl<7> vdd vss wl<124> / cell_PIM2
XI17968 bl<13> cbl<6> in1<110> in2<110> sl<13> vdd vss wl<110> / cell_PIM2
XI17967 bl<13> cbl<6> in1<109> in2<109> sl<13> vdd vss wl<109> / cell_PIM2
XI17966 bl<13> cbl<6> in1<108> in2<108> sl<13> vdd vss wl<108> / cell_PIM2
XI17965 bl<13> cbl<6> in1<107> in2<107> sl<13> vdd vss wl<107> / cell_PIM2
XI17964 bl<13> cbl<6> in1<106> in2<106> sl<13> vdd vss wl<106> / cell_PIM2
XI18618 bl<13> cbl<6> in1<28> in2<28> sl<13> vdd vss wl<28> / cell_PIM2
XI18617 bl<13> cbl<6> in1<27> in2<27> sl<13> vdd vss wl<27> / cell_PIM2
XI18616 bl<13> cbl<6> in1<26> in2<26> sl<13> vdd vss wl<26> / cell_PIM2
XI18615 bl<13> cbl<6> in1<25> in2<25> sl<13> vdd vss wl<25> / cell_PIM2
XI17312 bl<5> cbl<2> in1<124> in2<124> sl<5> vdd vss wl<124> / cell_PIM2
XI17311 bl<5> cbl<2> in1<123> in2<123> sl<5> vdd vss wl<123> / cell_PIM2
XI17310 bl<5> cbl<2> in1<122> in2<122> sl<5> vdd vss wl<122> / cell_PIM2
XI17309 bl<5> cbl<2> in1<121> in2<121> sl<5> vdd vss wl<121> / cell_PIM2
XI18610 bl<11> cbl<5> in1<25> in2<25> sl<11> vdd vss wl<25> / cell_PIM2
XI18609 bl<11> cbl<5> in1<26> in2<26> sl<11> vdd vss wl<26> / cell_PIM2
XI18608 bl<11> cbl<5> in1<27> in2<27> sl<11> vdd vss wl<27> / cell_PIM2
XI18607 bl<11> cbl<5> in1<28> in2<28> sl<11> vdd vss wl<28> / cell_PIM2
XI17958 bl<11> cbl<5> in1<106> in2<106> sl<11> vdd vss wl<106> / cell_PIM2
XI17957 bl<11> cbl<5> in1<107> in2<107> sl<11> vdd vss wl<107> / cell_PIM2
XI17956 bl<11> cbl<5> in1<108> in2<108> sl<11> vdd vss wl<108> / cell_PIM2
XI17955 bl<11> cbl<5> in1<109> in2<109> sl<11> vdd vss wl<109> / cell_PIM2
XI17954 bl<11> cbl<5> in1<110> in2<110> sl<11> vdd vss wl<110> / cell_PIM2
XI17308 bl<5> cbl<2> in1<120> in2<120> sl<5> vdd vss wl<120> / cell_PIM2
XI17302 bl<7> cbl<3> in1<127> in2<127> sl<7> vdd vss wl<127> / cell_PIM2
XI17301 bl<7> cbl<3> in1<126> in2<126> sl<7> vdd vss wl<126> / cell_PIM2
XI17300 bl<7> cbl<3> in1<125> in2<125> sl<7> vdd vss wl<125> / cell_PIM2
XI18602 bl<9> cbl<4> in1<28> in2<28> sl<9> vdd vss wl<28> / cell_PIM2
XI18601 bl<9> cbl<4> in1<27> in2<27> sl<9> vdd vss wl<27> / cell_PIM2
XI18600 bl<9> cbl<4> in1<26> in2<26> sl<9> vdd vss wl<26> / cell_PIM2
XI18599 bl<9> cbl<4> in1<25> in2<25> sl<9> vdd vss wl<25> / cell_PIM2
XI17296 bl<5> cbl<2> in1<127> in2<127> sl<5> vdd vss wl<127> / cell_PIM2
XI17295 bl<5> cbl<2> in1<126> in2<126> sl<5> vdd vss wl<126> / cell_PIM2
XI17294 bl<5> cbl<2> in1<125> in2<125> sl<5> vdd vss wl<125> / cell_PIM2
XI17948 bl<9> cbl<4> in1<110> in2<110> sl<9> vdd vss wl<110> / cell_PIM2
XI17947 bl<9> cbl<4> in1<109> in2<109> sl<9> vdd vss wl<109> / cell_PIM2
XI17946 bl<9> cbl<4> in1<108> in2<108> sl<9> vdd vss wl<108> / cell_PIM2
XI17945 bl<9> cbl<4> in1<107> in2<107> sl<9> vdd vss wl<107> / cell_PIM2
XI17944 bl<9> cbl<4> in1<106> in2<106> sl<9> vdd vss wl<106> / cell_PIM2
XI18594 bl<15> cbl<7> in1<29> in2<29> sl<15> vdd vss wl<29> / cell_PIM2
XI17289 bl<3> cbl<1> in1<0> in2<0> sl<3> vdd vss wl<0> / cell_PIM2
XI18593 bl<15> cbl<7> in1<30> in2<30> sl<15> vdd vss wl<30> / cell_PIM2
XI18592 bl<15> cbl<7> in1<31> in2<31> sl<15> vdd vss wl<31> / cell_PIM2
XI18591 bl<15> cbl<7> in1<32> in2<32> sl<15> vdd vss wl<32> / cell_PIM2
XI18590 bl<15> cbl<7> in1<33> in2<33> sl<15> vdd vss wl<33> / cell_PIM2
XI18584 bl<13> cbl<6> in1<33> in2<33> sl<13> vdd vss wl<33> / cell_PIM2
XI17938 bl<15> cbl<7> in1<111> in2<111> sl<15> vdd vss wl<111> / cell_PIM2
XI17937 bl<15> cbl<7> in1<112> in2<112> sl<15> vdd vss wl<112> / cell_PIM2
XI17936 bl<15> cbl<7> in1<113> in2<113> sl<15> vdd vss wl<113> / cell_PIM2
XI17935 bl<15> cbl<7> in1<114> in2<114> sl<15> vdd vss wl<114> / cell_PIM2
XI17934 bl<15> cbl<7> in1<115> in2<115> sl<15> vdd vss wl<115> / cell_PIM2
XI17284 bl<3> cbl<1> in1<2> in2<2> sl<3> vdd vss wl<2> / cell_PIM2
XI17283 bl<3> cbl<1> in1<3> in2<3> sl<3> vdd vss wl<3> / cell_PIM2
XI17282 bl<3> cbl<1> in1<4> in2<4> sl<3> vdd vss wl<4> / cell_PIM2
XI17281 bl<3> cbl<1> in1<1> in2<1> sl<3> vdd vss wl<1> / cell_PIM2
XI17280 bl<3> cbl<1> in1<9> in2<9> sl<3> vdd vss wl<9> / cell_PIM2
XI17279 bl<3> cbl<1> in1<8> in2<8> sl<3> vdd vss wl<8> / cell_PIM2
XI18583 bl<13> cbl<6> in1<32> in2<32> sl<13> vdd vss wl<32> / cell_PIM2
XI18582 bl<13> cbl<6> in1<31> in2<31> sl<13> vdd vss wl<31> / cell_PIM2
XI18581 bl<13> cbl<6> in1<30> in2<30> sl<13> vdd vss wl<30> / cell_PIM2
XI18580 bl<13> cbl<6> in1<29> in2<29> sl<13> vdd vss wl<29> / cell_PIM2
XI17278 bl<3> cbl<1> in1<7> in2<7> sl<3> vdd vss wl<7> / cell_PIM2
XI17277 bl<3> cbl<1> in1<6> in2<6> sl<3> vdd vss wl<6> / cell_PIM2
XI17276 bl<3> cbl<1> in1<5> in2<5> sl<3> vdd vss wl<5> / cell_PIM2
XI17928 bl<13> cbl<6> in1<115> in2<115> sl<13> vdd vss wl<115> / cell_PIM2
XI17927 bl<13> cbl<6> in1<114> in2<114> sl<13> vdd vss wl<114> / cell_PIM2
XI17926 bl<13> cbl<6> in1<113> in2<113> sl<13> vdd vss wl<113> / cell_PIM2
XI17925 bl<13> cbl<6> in1<112> in2<112> sl<13> vdd vss wl<112> / cell_PIM2
XI17924 bl<13> cbl<6> in1<111> in2<111> sl<13> vdd vss wl<111> / cell_PIM2
XI18574 bl<11> cbl<5> in1<29> in2<29> sl<11> vdd vss wl<29> / cell_PIM2
XI17270 bl<3> cbl<1> in1<14> in2<14> sl<3> vdd vss wl<14> / cell_PIM2
XI17269 bl<3> cbl<1> in1<13> in2<13> sl<3> vdd vss wl<13> / cell_PIM2
XI18573 bl<11> cbl<5> in1<30> in2<30> sl<11> vdd vss wl<30> / cell_PIM2
XI18572 bl<11> cbl<5> in1<31> in2<31> sl<11> vdd vss wl<31> / cell_PIM2
XI18571 bl<11> cbl<5> in1<32> in2<32> sl<11> vdd vss wl<32> / cell_PIM2
XI18570 bl<11> cbl<5> in1<33> in2<33> sl<11> vdd vss wl<33> / cell_PIM2
XI18564 bl<9> cbl<4> in1<33> in2<33> sl<9> vdd vss wl<33> / cell_PIM2
XI17918 bl<11> cbl<5> in1<111> in2<111> sl<11> vdd vss wl<111> / cell_PIM2
XI17917 bl<11> cbl<5> in1<112> in2<112> sl<11> vdd vss wl<112> / cell_PIM2
XI17916 bl<11> cbl<5> in1<113> in2<113> sl<11> vdd vss wl<113> / cell_PIM2
XI17915 bl<11> cbl<5> in1<114> in2<114> sl<11> vdd vss wl<114> / cell_PIM2
XI17914 bl<11> cbl<5> in1<115> in2<115> sl<11> vdd vss wl<115> / cell_PIM2
XI17268 bl<3> cbl<1> in1<12> in2<12> sl<3> vdd vss wl<12> / cell_PIM2
XI17267 bl<3> cbl<1> in1<11> in2<11> sl<3> vdd vss wl<11> / cell_PIM2
XI17266 bl<3> cbl<1> in1<10> in2<10> sl<3> vdd vss wl<10> / cell_PIM2
XI17260 bl<3> cbl<1> in1<19> in2<19> sl<3> vdd vss wl<19> / cell_PIM2
XI17259 bl<3> cbl<1> in1<18> in2<18> sl<3> vdd vss wl<18> / cell_PIM2
XI18563 bl<9> cbl<4> in1<32> in2<32> sl<9> vdd vss wl<32> / cell_PIM2
XI18562 bl<9> cbl<4> in1<31> in2<31> sl<9> vdd vss wl<31> / cell_PIM2
XI18561 bl<9> cbl<4> in1<30> in2<30> sl<9> vdd vss wl<30> / cell_PIM2
XI18560 bl<9> cbl<4> in1<29> in2<29> sl<9> vdd vss wl<29> / cell_PIM2
XI17258 bl<3> cbl<1> in1<17> in2<17> sl<3> vdd vss wl<17> / cell_PIM2
XI17257 bl<3> cbl<1> in1<16> in2<16> sl<3> vdd vss wl<16> / cell_PIM2
XI17256 bl<3> cbl<1> in1<15> in2<15> sl<3> vdd vss wl<15> / cell_PIM2
XI17908 bl<9> cbl<4> in1<115> in2<115> sl<9> vdd vss wl<115> / cell_PIM2
XI17907 bl<9> cbl<4> in1<114> in2<114> sl<9> vdd vss wl<114> / cell_PIM2
XI17906 bl<9> cbl<4> in1<113> in2<113> sl<9> vdd vss wl<113> / cell_PIM2
XI17905 bl<9> cbl<4> in1<112> in2<112> sl<9> vdd vss wl<112> / cell_PIM2
XI17904 bl<9> cbl<4> in1<111> in2<111> sl<9> vdd vss wl<111> / cell_PIM2
XI18554 bl<15> cbl<7> in1<34> in2<34> sl<15> vdd vss wl<34> / cell_PIM2
XI22954 bl<47> cbl<23> in1<61> in2<61> sl<47> vdd vss wl<61> / cell_PIM2
XI22953 bl<47> cbl<23> in1<62> in2<62> sl<47> vdd vss wl<62> / cell_PIM2
XI24142 bl<39> cbl<19> in1<26> in2<26> sl<39> vdd vss wl<26> / cell_PIM2
XI24143 bl<39> cbl<19> in1<25> in2<25> sl<39> vdd vss wl<25> / cell_PIM2
XI24792 bl<47> cbl<23> in1<5> in2<5> sl<47> vdd vss wl<5> / cell_PIM2
XI24791 bl<47> cbl<23> in1<6> in2<6> sl<47> vdd vss wl<6> / cell_PIM2
XI24790 bl<47> cbl<23> in1<7> in2<7> sl<47> vdd vss wl<7> / cell_PIM2
XI24793 bl<47> cbl<23> in1<3> in2<3> sl<47> vdd vss wl<3> / cell_PIM2
XI24784 bl<45> cbl<22> in1<3> in2<3> sl<45> vdd vss wl<3> / cell_PIM2
XI24136 bl<37> cbl<18> in1<24> in2<24> sl<37> vdd vss wl<24> / cell_PIM2
XI24135 bl<37> cbl<18> in1<23> in2<23> sl<37> vdd vss wl<23> / cell_PIM2
XI24134 bl<37> cbl<18> in1<22> in2<22> sl<37> vdd vss wl<22> / cell_PIM2
XI23488 bl<61> cbl<30> in1<47> in2<47> sl<61> vdd vss wl<47> / cell_PIM2
XI23487 bl<61> cbl<30> in1<46> in2<46> sl<61> vdd vss wl<46> / cell_PIM2
XI23486 bl<61> cbl<30> in1<50> in2<50> sl<61> vdd vss wl<50> / cell_PIM2
XI23485 bl<61> cbl<30> in1<49> in2<49> sl<61> vdd vss wl<49> / cell_PIM2
XI23484 bl<61> cbl<30> in1<48> in2<48> sl<61> vdd vss wl<48> / cell_PIM2
XI22952 bl<47> cbl<23> in1<63> in2<63> sl<47> vdd vss wl<63> / cell_PIM2
XI22951 bl<47> cbl<23> in1<64> in2<64> sl<47> vdd vss wl<64> / cell_PIM2
XI22313 bl<39> cbl<19> in1<81> in2<81> sl<39> vdd vss wl<81> / cell_PIM2
XI22946 bl<45> cbl<22> in1<62> in2<62> sl<45> vdd vss wl<62> / cell_PIM2
XI22945 bl<45> cbl<22> in1<61> in2<61> sl<45> vdd vss wl<61> / cell_PIM2
XI24132 bl<37> cbl<18> in1<25> in2<25> sl<37> vdd vss wl<25> / cell_PIM2
XI24133 bl<37> cbl<18> in1<26> in2<26> sl<37> vdd vss wl<26> / cell_PIM2
XI24782 bl<45> cbl<22> in1<7> in2<7> sl<45> vdd vss wl<7> / cell_PIM2
XI24781 bl<45> cbl<22> in1<6> in2<6> sl<45> vdd vss wl<6> / cell_PIM2
XI24780 bl<45> cbl<22> in1<5> in2<5> sl<45> vdd vss wl<5> / cell_PIM2
XI24783 bl<45> cbl<22> in1<4> in2<4> sl<45> vdd vss wl<4> / cell_PIM2
XI22944 bl<45> cbl<22> in1<64> in2<64> sl<45> vdd vss wl<64> / cell_PIM2
XI22943 bl<45> cbl<22> in1<63> in2<63> sl<45> vdd vss wl<63> / cell_PIM2
XI23478 bl<59> cbl<29> in1<46> in2<46> sl<59> vdd vss wl<46> / cell_PIM2
XI23477 bl<59> cbl<29> in1<47> in2<47> sl<59> vdd vss wl<47> / cell_PIM2
XI23476 bl<59> cbl<29> in1<48> in2<48> sl<59> vdd vss wl<48> / cell_PIM2
XI23475 bl<59> cbl<29> in1<49> in2<49> sl<59> vdd vss wl<49> / cell_PIM2
XI23474 bl<59> cbl<29> in1<50> in2<50> sl<59> vdd vss wl<50> / cell_PIM2
XI24126 bl<35> cbl<17> in1<22> in2<22> sl<35> vdd vss wl<22> / cell_PIM2
XI24125 bl<35> cbl<17> in1<23> in2<23> sl<35> vdd vss wl<23> / cell_PIM2
XI24124 bl<35> cbl<17> in1<24> in2<24> sl<35> vdd vss wl<24> / cell_PIM2
XI24774 bl<43> cbl<21> in1<4> in2<4> sl<43> vdd vss wl<4> / cell_PIM2
XI22303 bl<37> cbl<18> in1<82> in2<82> sl<37> vdd vss wl<82> / cell_PIM2
XI22938 bl<43> cbl<21> in1<61> in2<61> sl<43> vdd vss wl<61> / cell_PIM2
XI22937 bl<43> cbl<21> in1<62> in2<62> sl<43> vdd vss wl<62> / cell_PIM2
XI24122 bl<35> cbl<17> in1<26> in2<26> sl<35> vdd vss wl<26> / cell_PIM2
XI24123 bl<35> cbl<17> in1<25> in2<25> sl<35> vdd vss wl<25> / cell_PIM2
XI24772 bl<43> cbl<21> in1<5> in2<5> sl<43> vdd vss wl<5> / cell_PIM2
XI24771 bl<43> cbl<21> in1<6> in2<6> sl<43> vdd vss wl<6> / cell_PIM2
XI24770 bl<43> cbl<21> in1<7> in2<7> sl<43> vdd vss wl<7> / cell_PIM2
XI24773 bl<43> cbl<21> in1<3> in2<3> sl<43> vdd vss wl<3> / cell_PIM2
XI24764 bl<41> cbl<20> in1<4> in2<4> sl<41> vdd vss wl<4> / cell_PIM2
XI24116 bl<33> cbl<16> in1<24> in2<24> sl<33> vdd vss wl<24> / cell_PIM2
XI24115 bl<33> cbl<16> in1<23> in2<23> sl<33> vdd vss wl<23> / cell_PIM2
XI24114 bl<33> cbl<16> in1<22> in2<22> sl<33> vdd vss wl<22> / cell_PIM2
XI23468 bl<57> cbl<28> in1<46> in2<46> sl<57> vdd vss wl<46> / cell_PIM2
XI23467 bl<57> cbl<28> in1<47> in2<47> sl<57> vdd vss wl<47> / cell_PIM2
XI23466 bl<57> cbl<28> in1<48> in2<48> sl<57> vdd vss wl<48> / cell_PIM2
XI23465 bl<57> cbl<28> in1<49> in2<49> sl<57> vdd vss wl<49> / cell_PIM2
XI23464 bl<57> cbl<28> in1<50> in2<50> sl<57> vdd vss wl<50> / cell_PIM2
XI22936 bl<43> cbl<21> in1<63> in2<63> sl<43> vdd vss wl<63> / cell_PIM2
XI22935 bl<43> cbl<21> in1<64> in2<64> sl<43> vdd vss wl<64> / cell_PIM2
XI22298 bl<35> cbl<17> in1<80> in2<80> sl<35> vdd vss wl<80> / cell_PIM2
XI22930 bl<41> cbl<20> in1<61> in2<61> sl<41> vdd vss wl<61> / cell_PIM2
XI22929 bl<41> cbl<20> in1<62> in2<62> sl<41> vdd vss wl<62> / cell_PIM2
XI24112 bl<33> cbl<16> in1<25> in2<25> sl<33> vdd vss wl<25> / cell_PIM2
XI24113 bl<33> cbl<16> in1<26> in2<26> sl<33> vdd vss wl<26> / cell_PIM2
XI24762 bl<41> cbl<20> in1<5> in2<5> sl<41> vdd vss wl<5> / cell_PIM2
XI24761 bl<41> cbl<20> in1<6> in2<6> sl<41> vdd vss wl<6> / cell_PIM2
XI24760 bl<41> cbl<20> in1<7> in2<7> sl<41> vdd vss wl<7> / cell_PIM2
XI24763 bl<41> cbl<20> in1<3> in2<3> sl<41> vdd vss wl<3> / cell_PIM2
XI22288 bl<33> cbl<16> in1<83> in2<83> sl<33> vdd vss wl<83> / cell_PIM2
XI22928 bl<41> cbl<20> in1<63> in2<63> sl<41> vdd vss wl<63> / cell_PIM2
XI22927 bl<41> cbl<20> in1<64> in2<64> sl<41> vdd vss wl<64> / cell_PIM2
XI23458 bl<55> cbl<27> in1<46> in2<46> sl<55> vdd vss wl<46> / cell_PIM2
XI23457 bl<55> cbl<27> in1<47> in2<47> sl<55> vdd vss wl<47> / cell_PIM2
XI23456 bl<55> cbl<27> in1<48> in2<48> sl<55> vdd vss wl<48> / cell_PIM2
XI23455 bl<55> cbl<27> in1<49> in2<49> sl<55> vdd vss wl<49> / cell_PIM2
XI23454 bl<55> cbl<27> in1<50> in2<50> sl<55> vdd vss wl<50> / cell_PIM2
XI24106 bl<63> cbl<31> in1<27> in2<27> sl<63> vdd vss wl<27> / cell_PIM2
XI24105 bl<63> cbl<31> in1<28> in2<28> sl<63> vdd vss wl<28> / cell_PIM2
XI24104 bl<63> cbl<31> in1<29> in2<29> sl<63> vdd vss wl<29> / cell_PIM2
XI24754 bl<39> cbl<19> in1<4> in2<4> sl<39> vdd vss wl<4> / cell_PIM2
XI17250 bl<3> cbl<1> in1<24> in2<24> sl<3> vdd vss wl<24> / cell_PIM2
XI17249 bl<3> cbl<1> in1<23> in2<23> sl<3> vdd vss wl<23> / cell_PIM2
XI18553 bl<15> cbl<7> in1<35> in2<35> sl<15> vdd vss wl<35> / cell_PIM2
XI18552 bl<15> cbl<7> in1<36> in2<36> sl<15> vdd vss wl<36> / cell_PIM2
XI18551 bl<15> cbl<7> in1<37> in2<37> sl<15> vdd vss wl<37> / cell_PIM2
XI18550 bl<15> cbl<7> in1<38> in2<38> sl<15> vdd vss wl<38> / cell_PIM2
XI19202 bl<29> cbl<14> in1<105> in2<105> sl<29> vdd vss wl<105> / cell_PIM2
XI19201 bl<29> cbl<14> in1<104> in2<104> sl<29> vdd vss wl<104> / cell_PIM2
XI19200 bl<29> cbl<14> in1<107> in2<107> sl<29> vdd vss wl<107> / cell_PIM2
XI19199 bl<29> cbl<14> in1<106> in2<106> sl<29> vdd vss wl<106> / cell_PIM2
XI19834 bl<31> cbl<15> in1<65> in2<65> sl<31> vdd vss wl<65> / cell_PIM2
XI19833 bl<31> cbl<15> in1<66> in2<66> sl<31> vdd vss wl<66> / cell_PIM2
XI20372 bl<17> cbl<8> in1<28> in2<28> sl<17> vdd vss wl<28> / cell_PIM2
XI20371 bl<17> cbl<8> in1<27> in2<27> sl<17> vdd vss wl<27> / cell_PIM2
XI20370 bl<17> cbl<8> in1<31> in2<31> sl<17> vdd vss wl<31> / cell_PIM2
XI20369 bl<17> cbl<8> in1<30> in2<30> sl<17> vdd vss wl<30> / cell_PIM2
XI21023 bl<61> cbl<30> in1<126> in2<126> sl<61> vdd vss wl<126> / cell_PIM2
XI21022 bl<61> cbl<30> in1<125> in2<125> sl<61> vdd vss wl<125> / cell_PIM2
XI21021 bl<61> cbl<30> in1<124> in2<124> sl<61> vdd vss wl<124> / cell_PIM2
XI21020 bl<61> cbl<30> in1<123> in2<123> sl<61> vdd vss wl<123> / cell_PIM2
XI21672 bl<37> cbl<18> in1<100> in2<100> sl<37> vdd vss wl<100> / cell_PIM2
XI21671 bl<37> cbl<18> in1<99> in2<99> sl<37> vdd vss wl<99> / cell_PIM2
XI21670 bl<37> cbl<18> in1<103> in2<103> sl<37> vdd vss wl<103> / cell_PIM2
XI21669 bl<37> cbl<18> in1<102> in2<102> sl<37> vdd vss wl<102> / cell_PIM2
XI22322 bl<41> cbl<20> in1<80> in2<80> sl<41> vdd vss wl<80> / cell_PIM2
XI22321 bl<41> cbl<20> in1<81> in2<81> sl<41> vdd vss wl<81> / cell_PIM2
XI22320 bl<41> cbl<20> in1<82> in2<82> sl<41> vdd vss wl<82> / cell_PIM2
XI22319 bl<41> cbl<20> in1<83> in2<83> sl<41> vdd vss wl<83> / cell_PIM2
XI21668 bl<37> cbl<18> in1<101> in2<101> sl<37> vdd vss wl<101> / cell_PIM2
XI21014 bl<59> cbl<29> in1<127> in2<127> sl<59> vdd vss wl<127> / cell_PIM2
XI20368 bl<17> cbl<8> in1<29> in2<29> sl<17> vdd vss wl<29> / cell_PIM2
XI19832 bl<31> cbl<15> in1<67> in2<67> sl<31> vdd vss wl<67> / cell_PIM2
XI19831 bl<31> cbl<15> in1<68> in2<68> sl<31> vdd vss wl<68> / cell_PIM2
XI19830 bl<31> cbl<15> in1<69> in2<69> sl<31> vdd vss wl<69> / cell_PIM2
XI19194 bl<27> cbl<13> in1<104> in2<104> sl<27> vdd vss wl<104> / cell_PIM2
XI18544 bl<13> cbl<6> in1<38> in2<38> sl<13> vdd vss wl<38> / cell_PIM2
XI17898 bl<15> cbl<7> in1<116> in2<116> sl<15> vdd vss wl<116> / cell_PIM2
XI17897 bl<15> cbl<7> in1<117> in2<117> sl<15> vdd vss wl<117> / cell_PIM2
XI17896 bl<15> cbl<7> in1<118> in2<118> sl<15> vdd vss wl<118> / cell_PIM2
XI17895 bl<15> cbl<7> in1<119> in2<119> sl<15> vdd vss wl<119> / cell_PIM2
XI17248 bl<3> cbl<1> in1<22> in2<22> sl<3> vdd vss wl<22> / cell_PIM2
XI17247 bl<3> cbl<1> in1<21> in2<21> sl<3> vdd vss wl<21> / cell_PIM2
XI17246 bl<3> cbl<1> in1<20> in2<20> sl<3> vdd vss wl<20> / cell_PIM2
XI22314 bl<39> cbl<19> in1<80> in2<80> sl<39> vdd vss wl<80> / cell_PIM2
XI17240 bl<3> cbl<1> in1<28> in2<28> sl<3> vdd vss wl<28> / cell_PIM2
XI17239 bl<3> cbl<1> in1<27> in2<27> sl<3> vdd vss wl<27> / cell_PIM2
XI17890 bl<13> cbl<6> in1<119> in2<119> sl<13> vdd vss wl<119> / cell_PIM2
XI17889 bl<13> cbl<6> in1<118> in2<118> sl<13> vdd vss wl<118> / cell_PIM2
XI18543 bl<13> cbl<6> in1<37> in2<37> sl<13> vdd vss wl<37> / cell_PIM2
XI18542 bl<13> cbl<6> in1<36> in2<36> sl<13> vdd vss wl<36> / cell_PIM2
XI18541 bl<13> cbl<6> in1<35> in2<35> sl<13> vdd vss wl<35> / cell_PIM2
XI18540 bl<13> cbl<6> in1<34> in2<34> sl<13> vdd vss wl<34> / cell_PIM2
XI19192 bl<27> cbl<13> in1<106> in2<106> sl<27> vdd vss wl<106> / cell_PIM2
XI19191 bl<27> cbl<13> in1<107> in2<107> sl<27> vdd vss wl<107> / cell_PIM2
XI19193 bl<27> cbl<13> in1<105> in2<105> sl<27> vdd vss wl<105> / cell_PIM2
XI20362 bl<31> cbl<15> in1<32> in2<32> sl<31> vdd vss wl<32> / cell_PIM2
XI20361 bl<31> cbl<15> in1<33> in2<33> sl<31> vdd vss wl<33> / cell_PIM2
XI20360 bl<31> cbl<15> in1<34> in2<34> sl<31> vdd vss wl<34> / cell_PIM2
XI20359 bl<31> cbl<15> in1<35> in2<35> sl<31> vdd vss wl<35> / cell_PIM2
XI21013 bl<59> cbl<29> in1<126> in2<126> sl<59> vdd vss wl<126> / cell_PIM2
XI21012 bl<59> cbl<29> in1<125> in2<125> sl<59> vdd vss wl<125> / cell_PIM2
XI21011 bl<59> cbl<29> in1<123> in2<123> sl<59> vdd vss wl<123> / cell_PIM2
XI21010 bl<59> cbl<29> in1<124> in2<124> sl<59> vdd vss wl<124> / cell_PIM2
XI21662 bl<35> cbl<17> in1<99> in2<99> sl<35> vdd vss wl<99> / cell_PIM2
XI21661 bl<35> cbl<17> in1<100> in2<100> sl<35> vdd vss wl<100> / cell_PIM2
XI21660 bl<35> cbl<17> in1<101> in2<101> sl<35> vdd vss wl<101> / cell_PIM2
XI21659 bl<35> cbl<17> in1<102> in2<102> sl<35> vdd vss wl<102> / cell_PIM2
XI22312 bl<39> cbl<19> in1<82> in2<82> sl<39> vdd vss wl<82> / cell_PIM2
XI22311 bl<39> cbl<19> in1<83> in2<83> sl<39> vdd vss wl<83> / cell_PIM2
XI17238 bl<3> cbl<1> in1<26> in2<26> sl<3> vdd vss wl<26> / cell_PIM2
XI17237 bl<3> cbl<1> in1<25> in2<25> sl<3> vdd vss wl<25> / cell_PIM2
XI17888 bl<13> cbl<6> in1<117> in2<117> sl<13> vdd vss wl<117> / cell_PIM2
XI17887 bl<13> cbl<6> in1<116> in2<116> sl<13> vdd vss wl<116> / cell_PIM2
XI18534 bl<11> cbl<5> in1<34> in2<34> sl<11> vdd vss wl<34> / cell_PIM2
XI19186 bl<25> cbl<12> in1<104> in2<104> sl<25> vdd vss wl<104> / cell_PIM2
XI19185 bl<25> cbl<12> in1<105> in2<105> sl<25> vdd vss wl<105> / cell_PIM2
XI19184 bl<25> cbl<12> in1<106> in2<106> sl<25> vdd vss wl<106> / cell_PIM2
XI19824 bl<29> cbl<14> in1<67> in2<67> sl<29> vdd vss wl<67> / cell_PIM2
XI19823 bl<29> cbl<14> in1<66> in2<66> sl<29> vdd vss wl<66> / cell_PIM2
XI19822 bl<29> cbl<14> in1<65> in2<65> sl<29> vdd vss wl<65> / cell_PIM2
XI19821 bl<29> cbl<14> in1<69> in2<69> sl<29> vdd vss wl<69> / cell_PIM2
XI20358 bl<31> cbl<15> in1<36> in2<36> sl<31> vdd vss wl<36> / cell_PIM2
XI21004 bl<57> cbl<28> in1<127> in2<127> sl<57> vdd vss wl<127> / cell_PIM2
XI21658 bl<35> cbl<17> in1<103> in2<103> sl<35> vdd vss wl<103> / cell_PIM2
XI22306 bl<37> cbl<18> in1<81> in2<81> sl<37> vdd vss wl<81> / cell_PIM2
XI22305 bl<37> cbl<18> in1<80> in2<80> sl<37> vdd vss wl<80> / cell_PIM2
XI22304 bl<37> cbl<18> in1<83> in2<83> sl<37> vdd vss wl<83> / cell_PIM2
XI17232 bl<3> cbl<1> in1<33> in2<33> sl<3> vdd vss wl<33> / cell_PIM2
XI17231 bl<3> cbl<1> in1<32> in2<32> sl<3> vdd vss wl<32> / cell_PIM2
XI17230 bl<3> cbl<1> in1<31> in2<31> sl<3> vdd vss wl<31> / cell_PIM2
XI17229 bl<3> cbl<1> in1<30> in2<30> sl<3> vdd vss wl<30> / cell_PIM2
XI17882 bl<11> cbl<5> in1<116> in2<116> sl<11> vdd vss wl<116> / cell_PIM2
XI17881 bl<11> cbl<5> in1<117> in2<117> sl<11> vdd vss wl<117> / cell_PIM2
XI17880 bl<11> cbl<5> in1<118> in2<118> sl<11> vdd vss wl<118> / cell_PIM2
XI17879 bl<11> cbl<5> in1<119> in2<119> sl<11> vdd vss wl<119> / cell_PIM2
XI18533 bl<11> cbl<5> in1<35> in2<35> sl<11> vdd vss wl<35> / cell_PIM2
XI18532 bl<11> cbl<5> in1<36> in2<36> sl<11> vdd vss wl<36> / cell_PIM2
XI18531 bl<11> cbl<5> in1<37> in2<37> sl<11> vdd vss wl<37> / cell_PIM2
XI18530 bl<11> cbl<5> in1<38> in2<38> sl<11> vdd vss wl<38> / cell_PIM2
XI19183 bl<25> cbl<12> in1<107> in2<107> sl<25> vdd vss wl<107> / cell_PIM2
XI19820 bl<29> cbl<14> in1<68> in2<68> sl<29> vdd vss wl<68> / cell_PIM2
XI20352 bl<29> cbl<14> in1<33> in2<33> sl<29> vdd vss wl<33> / cell_PIM2
XI20351 bl<29> cbl<14> in1<32> in2<32> sl<29> vdd vss wl<32> / cell_PIM2
XI20350 bl<29> cbl<14> in1<36> in2<36> sl<29> vdd vss wl<36> / cell_PIM2
XI20349 bl<29> cbl<14> in1<35> in2<35> sl<29> vdd vss wl<35> / cell_PIM2
XI21003 bl<57> cbl<28> in1<126> in2<126> sl<57> vdd vss wl<126> / cell_PIM2
XI21002 bl<57> cbl<28> in1<125> in2<125> sl<57> vdd vss wl<125> / cell_PIM2
XI21001 bl<57> cbl<28> in1<123> in2<123> sl<57> vdd vss wl<123> / cell_PIM2
XI21000 bl<57> cbl<28> in1<124> in2<124> sl<57> vdd vss wl<124> / cell_PIM2
XI21652 bl<33> cbl<16> in1<100> in2<100> sl<33> vdd vss wl<100> / cell_PIM2
XI21651 bl<33> cbl<16> in1<99> in2<99> sl<33> vdd vss wl<99> / cell_PIM2
XI21650 bl<33> cbl<16> in1<103> in2<103> sl<33> vdd vss wl<103> / cell_PIM2
XI21649 bl<33> cbl<16> in1<102> in2<102> sl<33> vdd vss wl<102> / cell_PIM2
XI22297 bl<35> cbl<17> in1<81> in2<81> sl<35> vdd vss wl<81> / cell_PIM2
XI22296 bl<35> cbl<17> in1<82> in2<82> sl<35> vdd vss wl<82> / cell_PIM2
XI22295 bl<35> cbl<17> in1<83> in2<83> sl<35> vdd vss wl<83> / cell_PIM2
XI21648 bl<33> cbl<16> in1<101> in2<101> sl<33> vdd vss wl<101> / cell_PIM2
XI20994 bl<55> cbl<27> in1<127> in2<127> sl<55> vdd vss wl<127> / cell_PIM2
XI20348 bl<29> cbl<14> in1<34> in2<34> sl<29> vdd vss wl<34> / cell_PIM2
XI19814 bl<27> cbl<13> in1<65> in2<65> sl<27> vdd vss wl<65> / cell_PIM2
XI19813 bl<27> cbl<13> in1<66> in2<66> sl<27> vdd vss wl<66> / cell_PIM2
XI19178 bl<23> cbl<11> in1<104> in2<104> sl<23> vdd vss wl<104> / cell_PIM2
XI19177 bl<23> cbl<11> in1<105> in2<105> sl<23> vdd vss wl<105> / cell_PIM2
XI19176 bl<23> cbl<11> in1<106> in2<106> sl<23> vdd vss wl<106> / cell_PIM2
XI19175 bl<23> cbl<11> in1<107> in2<107> sl<23> vdd vss wl<107> / cell_PIM2
XI18524 bl<9> cbl<4> in1<38> in2<38> sl<9> vdd vss wl<38> / cell_PIM2
XI17874 bl<9> cbl<4> in1<119> in2<119> sl<9> vdd vss wl<119> / cell_PIM2
XI17228 bl<3> cbl<1> in1<29> in2<29> sl<3> vdd vss wl<29> / cell_PIM2
XI17222 bl<3> cbl<1> in1<38> in2<38> sl<3> vdd vss wl<38> / cell_PIM2
XI17221 bl<3> cbl<1> in1<37> in2<37> sl<3> vdd vss wl<37> / cell_PIM2
XI17220 bl<3> cbl<1> in1<36> in2<36> sl<3> vdd vss wl<36> / cell_PIM2
XI17219 bl<3> cbl<1> in1<35> in2<35> sl<3> vdd vss wl<35> / cell_PIM2
XI17873 bl<9> cbl<4> in1<118> in2<118> sl<9> vdd vss wl<118> / cell_PIM2
XI17872 bl<9> cbl<4> in1<117> in2<117> sl<9> vdd vss wl<117> / cell_PIM2
XI17871 bl<9> cbl<4> in1<116> in2<116> sl<9> vdd vss wl<116> / cell_PIM2
XI18523 bl<9> cbl<4> in1<37> in2<37> sl<9> vdd vss wl<37> / cell_PIM2
XI18522 bl<9> cbl<4> in1<36> in2<36> sl<9> vdd vss wl<36> / cell_PIM2
XI18521 bl<9> cbl<4> in1<35> in2<35> sl<9> vdd vss wl<35> / cell_PIM2
XI18520 bl<9> cbl<4> in1<34> in2<34> sl<9> vdd vss wl<34> / cell_PIM2
XI19170 bl<21> cbl<10> in1<105> in2<105> sl<21> vdd vss wl<105> / cell_PIM2
XI19169 bl<21> cbl<10> in1<104> in2<104> sl<21> vdd vss wl<104> / cell_PIM2
XI19812 bl<27> cbl<13> in1<67> in2<67> sl<27> vdd vss wl<67> / cell_PIM2
XI19811 bl<27> cbl<13> in1<68> in2<68> sl<27> vdd vss wl<68> / cell_PIM2
XI19810 bl<27> cbl<13> in1<69> in2<69> sl<27> vdd vss wl<69> / cell_PIM2
XI20342 bl<27> cbl<13> in1<32> in2<32> sl<27> vdd vss wl<32> / cell_PIM2
XI20341 bl<27> cbl<13> in1<33> in2<33> sl<27> vdd vss wl<33> / cell_PIM2
XI20340 bl<27> cbl<13> in1<34> in2<34> sl<27> vdd vss wl<34> / cell_PIM2
XI20339 bl<27> cbl<13> in1<35> in2<35> sl<27> vdd vss wl<35> / cell_PIM2
XI20993 bl<55> cbl<27> in1<126> in2<126> sl<55> vdd vss wl<126> / cell_PIM2
XI20992 bl<55> cbl<27> in1<125> in2<125> sl<55> vdd vss wl<125> / cell_PIM2
XI20991 bl<55> cbl<27> in1<123> in2<123> sl<55> vdd vss wl<123> / cell_PIM2
XI20990 bl<55> cbl<27> in1<124> in2<124> sl<55> vdd vss wl<124> / cell_PIM2
XI21642 bl<63> cbl<31> in1<104> in2<104> sl<63> vdd vss wl<104> / cell_PIM2
XI21641 bl<63> cbl<31> in1<105> in2<105> sl<63> vdd vss wl<105> / cell_PIM2
XI21640 bl<63> cbl<31> in1<106> in2<106> sl<63> vdd vss wl<106> / cell_PIM2
XI21639 bl<63> cbl<31> in1<107> in2<107> sl<63> vdd vss wl<107> / cell_PIM2
XI22290 bl<33> cbl<16> in1<81> in2<81> sl<33> vdd vss wl<81> / cell_PIM2
XI22289 bl<33> cbl<16> in1<80> in2<80> sl<33> vdd vss wl<80> / cell_PIM2
XI17218 bl<3> cbl<1> in1<34> in2<34> sl<3> vdd vss wl<34> / cell_PIM2
XI17866 bl<15> cbl<7> in1<120> in2<120> sl<15> vdd vss wl<120> / cell_PIM2
XI17865 bl<15> cbl<7> in1<121> in2<121> sl<15> vdd vss wl<121> / cell_PIM2
XI17864 bl<15> cbl<7> in1<122> in2<122> sl<15> vdd vss wl<122> / cell_PIM2
XI18514 bl<15> cbl<7> in1<39> in2<39> sl<15> vdd vss wl<39> / cell_PIM2
XI19167 bl<21> cbl<10> in1<106> in2<106> sl<21> vdd vss wl<106> / cell_PIM2
XI19168 bl<21> cbl<10> in1<107> in2<107> sl<21> vdd vss wl<107> / cell_PIM2
XI20338 bl<27> cbl<13> in1<36> in2<36> sl<27> vdd vss wl<36> / cell_PIM2
XI20984 bl<53> cbl<26> in1<127> in2<127> sl<53> vdd vss wl<127> / cell_PIM2
XI21634 bl<61> cbl<30> in1<105> in2<105> sl<61> vdd vss wl<105> / cell_PIM2
XI22287 bl<33> cbl<16> in1<82> in2<82> sl<33> vdd vss wl<82> / cell_PIM2
XI22922 bl<39> cbl<19> in1<61> in2<61> sl<39> vdd vss wl<61> / cell_PIM2
XI22921 bl<39> cbl<19> in1<62> in2<62> sl<39> vdd vss wl<62> / cell_PIM2
XI24102 bl<63> cbl<31> in1<31> in2<31> sl<63> vdd vss wl<31> / cell_PIM2
XI24103 bl<63> cbl<31> in1<30> in2<30> sl<63> vdd vss wl<30> / cell_PIM2
XI24752 bl<39> cbl<19> in1<5> in2<5> sl<39> vdd vss wl<5> / cell_PIM2
XI24751 bl<39> cbl<19> in1<6> in2<6> sl<39> vdd vss wl<6> / cell_PIM2
XI24750 bl<39> cbl<19> in1<7> in2<7> sl<39> vdd vss wl<7> / cell_PIM2
XI24753 bl<39> cbl<19> in1<3> in2<3> sl<39> vdd vss wl<3> / cell_PIM2
XI24744 bl<37> cbl<18> in1<3> in2<3> sl<37> vdd vss wl<3> / cell_PIM2
XI24096 bl<61> cbl<30> in1<28> in2<28> sl<61> vdd vss wl<28> / cell_PIM2
XI24095 bl<61> cbl<30> in1<27> in2<27> sl<61> vdd vss wl<27> / cell_PIM2
XI24094 bl<61> cbl<30> in1<31> in2<31> sl<61> vdd vss wl<31> / cell_PIM2
XI23448 bl<53> cbl<26> in1<47> in2<47> sl<53> vdd vss wl<47> / cell_PIM2
XI23447 bl<53> cbl<26> in1<46> in2<46> sl<53> vdd vss wl<46> / cell_PIM2
XI23446 bl<53> cbl<26> in1<50> in2<50> sl<53> vdd vss wl<50> / cell_PIM2
XI23445 bl<53> cbl<26> in1<49> in2<49> sl<53> vdd vss wl<49> / cell_PIM2
XI23444 bl<53> cbl<26> in1<48> in2<48> sl<53> vdd vss wl<48> / cell_PIM2
XI22920 bl<39> cbl<19> in1<63> in2<63> sl<39> vdd vss wl<63> / cell_PIM2
XI22919 bl<39> cbl<19> in1<64> in2<64> sl<39> vdd vss wl<64> / cell_PIM2
XI22278 bl<63> cbl<31> in1<88> in2<88> sl<63> vdd vss wl<88> / cell_PIM2
XI22914 bl<37> cbl<18> in1<62> in2<62> sl<37> vdd vss wl<62> / cell_PIM2
XI22913 bl<37> cbl<18> in1<61> in2<61> sl<37> vdd vss wl<61> / cell_PIM2
XI24092 bl<61> cbl<30> in1<29> in2<29> sl<61> vdd vss wl<29> / cell_PIM2
XI24093 bl<61> cbl<30> in1<30> in2<30> sl<61> vdd vss wl<30> / cell_PIM2
XI24742 bl<37> cbl<18> in1<7> in2<7> sl<37> vdd vss wl<7> / cell_PIM2
XI24741 bl<37> cbl<18> in1<6> in2<6> sl<37> vdd vss wl<6> / cell_PIM2
XI24740 bl<37> cbl<18> in1<5> in2<5> sl<37> vdd vss wl<5> / cell_PIM2
XI24743 bl<37> cbl<18> in1<4> in2<4> sl<37> vdd vss wl<4> / cell_PIM2
XI22268 bl<61> cbl<30> in1<87> in2<87> sl<61> vdd vss wl<87> / cell_PIM2
XI22912 bl<37> cbl<18> in1<64> in2<64> sl<37> vdd vss wl<64> / cell_PIM2
XI22911 bl<37> cbl<18> in1<63> in2<63> sl<37> vdd vss wl<63> / cell_PIM2
XI23438 bl<51> cbl<25> in1<46> in2<46> sl<51> vdd vss wl<46> / cell_PIM2
XI23437 bl<51> cbl<25> in1<47> in2<47> sl<51> vdd vss wl<47> / cell_PIM2
XI23436 bl<51> cbl<25> in1<48> in2<48> sl<51> vdd vss wl<48> / cell_PIM2
XI23435 bl<51> cbl<25> in1<49> in2<49> sl<51> vdd vss wl<49> / cell_PIM2
XI23434 bl<51> cbl<25> in1<50> in2<50> sl<51> vdd vss wl<50> / cell_PIM2
XI24086 bl<59> cbl<29> in1<27> in2<27> sl<59> vdd vss wl<27> / cell_PIM2
XI24085 bl<59> cbl<29> in1<28> in2<28> sl<59> vdd vss wl<28> / cell_PIM2
XI24084 bl<59> cbl<29> in1<29> in2<29> sl<59> vdd vss wl<29> / cell_PIM2
XI24734 bl<35> cbl<17> in1<4> in2<4> sl<35> vdd vss wl<4> / cell_PIM2
XI17212 bl<3> cbl<1> in1<43> in2<43> sl<3> vdd vss wl<43> / cell_PIM2
XI17211 bl<3> cbl<1> in1<42> in2<42> sl<3> vdd vss wl<42> / cell_PIM2
XI17210 bl<3> cbl<1> in1<41> in2<41> sl<3> vdd vss wl<41> / cell_PIM2
XI17209 bl<3> cbl<1> in1<40> in2<40> sl<3> vdd vss wl<40> / cell_PIM2
XI17863 bl<15> cbl<7> in1<123> in2<123> sl<15> vdd vss wl<123> / cell_PIM2
XI17862 bl<15> cbl<7> in1<124> in2<124> sl<15> vdd vss wl<124> / cell_PIM2
XI18513 bl<15> cbl<7> in1<40> in2<40> sl<15> vdd vss wl<40> / cell_PIM2
XI18512 bl<15> cbl<7> in1<41> in2<41> sl<15> vdd vss wl<41> / cell_PIM2
XI18511 bl<15> cbl<7> in1<42> in2<42> sl<15> vdd vss wl<42> / cell_PIM2
XI18510 bl<15> cbl<7> in1<43> in2<43> sl<15> vdd vss wl<43> / cell_PIM2
XI19162 bl<19> cbl<9> in1<104> in2<104> sl<19> vdd vss wl<104> / cell_PIM2
XI19161 bl<19> cbl<9> in1<105> in2<105> sl<19> vdd vss wl<105> / cell_PIM2
XI19160 bl<19> cbl<9> in1<106> in2<106> sl<19> vdd vss wl<106> / cell_PIM2
XI19159 bl<19> cbl<9> in1<107> in2<107> sl<19> vdd vss wl<107> / cell_PIM2
XI19804 bl<25> cbl<12> in1<65> in2<65> sl<25> vdd vss wl<65> / cell_PIM2
XI19803 bl<25> cbl<12> in1<66> in2<66> sl<25> vdd vss wl<66> / cell_PIM2
XI19802 bl<25> cbl<12> in1<67> in2<67> sl<25> vdd vss wl<67> / cell_PIM2
XI19801 bl<25> cbl<12> in1<68> in2<68> sl<25> vdd vss wl<68> / cell_PIM2
XI20332 bl<25> cbl<12> in1<32> in2<32> sl<25> vdd vss wl<32> / cell_PIM2
XI20331 bl<25> cbl<12> in1<33> in2<33> sl<25> vdd vss wl<33> / cell_PIM2
XI20330 bl<25> cbl<12> in1<34> in2<34> sl<25> vdd vss wl<34> / cell_PIM2
XI20329 bl<25> cbl<12> in1<35> in2<35> sl<25> vdd vss wl<35> / cell_PIM2
XI20983 bl<53> cbl<26> in1<126> in2<126> sl<53> vdd vss wl<126> / cell_PIM2
XI20982 bl<53> cbl<26> in1<125> in2<125> sl<53> vdd vss wl<125> / cell_PIM2
XI20981 bl<53> cbl<26> in1<124> in2<124> sl<53> vdd vss wl<124> / cell_PIM2
XI20980 bl<53> cbl<26> in1<123> in2<123> sl<53> vdd vss wl<123> / cell_PIM2
XI21632 bl<61> cbl<30> in1<107> in2<107> sl<61> vdd vss wl<107> / cell_PIM2
XI21631 bl<61> cbl<30> in1<106> in2<106> sl<61> vdd vss wl<106> / cell_PIM2
XI21633 bl<61> cbl<30> in1<104> in2<104> sl<61> vdd vss wl<104> / cell_PIM2
XI22282 bl<63> cbl<31> in1<84> in2<84> sl<63> vdd vss wl<84> / cell_PIM2
XI22281 bl<63> cbl<31> in1<85> in2<85> sl<63> vdd vss wl<85> / cell_PIM2
XI22280 bl<63> cbl<31> in1<86> in2<86> sl<63> vdd vss wl<86> / cell_PIM2
XI22279 bl<63> cbl<31> in1<87> in2<87> sl<63> vdd vss wl<87> / cell_PIM2
XI21626 bl<59> cbl<29> in1<104> in2<104> sl<59> vdd vss wl<104> / cell_PIM2
XI21625 bl<59> cbl<29> in1<105> in2<105> sl<59> vdd vss wl<105> / cell_PIM2
XI21624 bl<59> cbl<29> in1<106> in2<106> sl<59> vdd vss wl<106> / cell_PIM2
XI20974 bl<51> cbl<25> in1<127> in2<127> sl<51> vdd vss wl<127> / cell_PIM2
XI20328 bl<25> cbl<12> in1<36> in2<36> sl<25> vdd vss wl<36> / cell_PIM2
XI19800 bl<25> cbl<12> in1<69> in2<69> sl<25> vdd vss wl<69> / cell_PIM2
XI19154 bl<17> cbl<8> in1<105> in2<105> sl<17> vdd vss wl<105> / cell_PIM2
XI18504 bl<13> cbl<6> in1<43> in2<43> sl<13> vdd vss wl<43> / cell_PIM2
XI17856 bl<13> cbl<6> in1<124> in2<124> sl<13> vdd vss wl<124> / cell_PIM2
XI17855 bl<13> cbl<6> in1<123> in2<123> sl<13> vdd vss wl<123> / cell_PIM2
XI17854 bl<13> cbl<6> in1<122> in2<122> sl<13> vdd vss wl<122> / cell_PIM2
XI17208 bl<3> cbl<1> in1<39> in2<39> sl<3> vdd vss wl<39> / cell_PIM2
XI17202 bl<3> cbl<1> in1<47> in2<47> sl<3> vdd vss wl<47> / cell_PIM2
XI17201 bl<3> cbl<1> in1<46> in2<46> sl<3> vdd vss wl<46> / cell_PIM2
XI17200 bl<3> cbl<1> in1<45> in2<45> sl<3> vdd vss wl<45> / cell_PIM2
XI17199 bl<3> cbl<1> in1<44> in2<44> sl<3> vdd vss wl<44> / cell_PIM2
XI17853 bl<13> cbl<6> in1<121> in2<121> sl<13> vdd vss wl<121> / cell_PIM2
XI17852 bl<13> cbl<6> in1<120> in2<120> sl<13> vdd vss wl<120> / cell_PIM2
XI18503 bl<13> cbl<6> in1<42> in2<42> sl<13> vdd vss wl<42> / cell_PIM2
XI18502 bl<13> cbl<6> in1<41> in2<41> sl<13> vdd vss wl<41> / cell_PIM2
XI18501 bl<13> cbl<6> in1<40> in2<40> sl<13> vdd vss wl<40> / cell_PIM2
XI18500 bl<13> cbl<6> in1<39> in2<39> sl<13> vdd vss wl<39> / cell_PIM2
XI19152 bl<17> cbl<8> in1<107> in2<107> sl<17> vdd vss wl<107> / cell_PIM2
XI19151 bl<17> cbl<8> in1<106> in2<106> sl<17> vdd vss wl<106> / cell_PIM2
XI19153 bl<17> cbl<8> in1<104> in2<104> sl<17> vdd vss wl<104> / cell_PIM2
XI19794 bl<23> cbl<11> in1<65> in2<65> sl<23> vdd vss wl<65> / cell_PIM2
XI19793 bl<23> cbl<11> in1<66> in2<66> sl<23> vdd vss wl<66> / cell_PIM2
XI20322 bl<23> cbl<11> in1<32> in2<32> sl<23> vdd vss wl<32> / cell_PIM2
XI20321 bl<23> cbl<11> in1<33> in2<33> sl<23> vdd vss wl<33> / cell_PIM2
XI20320 bl<23> cbl<11> in1<34> in2<34> sl<23> vdd vss wl<34> / cell_PIM2
XI20319 bl<23> cbl<11> in1<35> in2<35> sl<23> vdd vss wl<35> / cell_PIM2
XI20973 bl<51> cbl<25> in1<126> in2<126> sl<51> vdd vss wl<126> / cell_PIM2
XI20972 bl<51> cbl<25> in1<125> in2<125> sl<51> vdd vss wl<125> / cell_PIM2
XI20971 bl<51> cbl<25> in1<123> in2<123> sl<51> vdd vss wl<123> / cell_PIM2
XI20970 bl<51> cbl<25> in1<124> in2<124> sl<51> vdd vss wl<124> / cell_PIM2
XI21623 bl<59> cbl<29> in1<107> in2<107> sl<59> vdd vss wl<107> / cell_PIM2
XI22272 bl<61> cbl<30> in1<86> in2<86> sl<61> vdd vss wl<86> / cell_PIM2
XI22271 bl<61> cbl<30> in1<85> in2<85> sl<61> vdd vss wl<85> / cell_PIM2
XI22270 bl<61> cbl<30> in1<84> in2<84> sl<61> vdd vss wl<84> / cell_PIM2
XI22269 bl<61> cbl<30> in1<88> in2<88> sl<61> vdd vss wl<88> / cell_PIM2
XI17194 bl<3> cbl<1> in1<52> in2<52> sl<3> vdd vss wl<52> / cell_PIM2
XI17846 bl<11> cbl<5> in1<120> in2<120> sl<11> vdd vss wl<120> / cell_PIM2
XI17845 bl<11> cbl<5> in1<121> in2<121> sl<11> vdd vss wl<121> / cell_PIM2
XI17844 bl<11> cbl<5> in1<122> in2<122> sl<11> vdd vss wl<122> / cell_PIM2
XI18494 bl<11> cbl<5> in1<39> in2<39> sl<11> vdd vss wl<39> / cell_PIM2
XI19146 bl<31> cbl<15> in1<108> in2<108> sl<31> vdd vss wl<108> / cell_PIM2
XI19145 bl<31> cbl<15> in1<109> in2<109> sl<31> vdd vss wl<109> / cell_PIM2
XI19144 bl<31> cbl<15> in1<110> in2<110> sl<31> vdd vss wl<110> / cell_PIM2
XI19792 bl<23> cbl<11> in1<67> in2<67> sl<23> vdd vss wl<67> / cell_PIM2
XI19791 bl<23> cbl<11> in1<68> in2<68> sl<23> vdd vss wl<68> / cell_PIM2
XI19790 bl<23> cbl<11> in1<69> in2<69> sl<23> vdd vss wl<69> / cell_PIM2
XI20318 bl<23> cbl<11> in1<36> in2<36> sl<23> vdd vss wl<36> / cell_PIM2
XI20964 bl<49> cbl<24> in1<127> in2<127> sl<49> vdd vss wl<127> / cell_PIM2
XI21617 bl<57> cbl<28> in1<105> in2<105> sl<57> vdd vss wl<105> / cell_PIM2
XI21616 bl<57> cbl<28> in1<106> in2<106> sl<57> vdd vss wl<106> / cell_PIM2
XI21615 bl<57> cbl<28> in1<107> in2<107> sl<57> vdd vss wl<107> / cell_PIM2
XI21618 bl<57> cbl<28> in1<104> in2<104> sl<57> vdd vss wl<104> / cell_PIM2
XI22906 bl<35> cbl<17> in1<61> in2<61> sl<35> vdd vss wl<61> / cell_PIM2
XI22905 bl<35> cbl<17> in1<62> in2<62> sl<35> vdd vss wl<62> / cell_PIM2
XI24082 bl<59> cbl<29> in1<31> in2<31> sl<59> vdd vss wl<31> / cell_PIM2
XI24083 bl<59> cbl<29> in1<30> in2<30> sl<59> vdd vss wl<30> / cell_PIM2
XI24732 bl<35> cbl<17> in1<5> in2<5> sl<35> vdd vss wl<5> / cell_PIM2
XI24731 bl<35> cbl<17> in1<6> in2<6> sl<35> vdd vss wl<6> / cell_PIM2
XI24730 bl<35> cbl<17> in1<7> in2<7> sl<35> vdd vss wl<7> / cell_PIM2
XI24733 bl<35> cbl<17> in1<3> in2<3> sl<35> vdd vss wl<3> / cell_PIM2
XI22258 bl<59> cbl<29> in1<88> in2<88> sl<59> vdd vss wl<88> / cell_PIM2
XI22903 bl<35> cbl<17> in1<64> in2<64> sl<35> vdd vss wl<64> / cell_PIM2
XI22904 bl<35> cbl<17> in1<63> in2<63> sl<35> vdd vss wl<63> / cell_PIM2
XI23424 bl<49> cbl<24> in1<48> in2<48> sl<49> vdd vss wl<48> / cell_PIM2
XI23425 bl<49> cbl<24> in1<49> in2<49> sl<49> vdd vss wl<49> / cell_PIM2
XI23426 bl<49> cbl<24> in1<50> in2<50> sl<49> vdd vss wl<50> / cell_PIM2
XI23427 bl<49> cbl<24> in1<46> in2<46> sl<49> vdd vss wl<46> / cell_PIM2
XI23428 bl<49> cbl<24> in1<47> in2<47> sl<49> vdd vss wl<47> / cell_PIM2
XI24074 bl<57> cbl<28> in1<29> in2<29> sl<57> vdd vss wl<29> / cell_PIM2
XI24075 bl<57> cbl<28> in1<28> in2<28> sl<57> vdd vss wl<28> / cell_PIM2
XI24076 bl<57> cbl<28> in1<27> in2<27> sl<57> vdd vss wl<27> / cell_PIM2
XI24724 bl<33> cbl<16> in1<3> in2<3> sl<33> vdd vss wl<3> / cell_PIM2
XI17193 bl<3> cbl<1> in1<51> in2<51> sl<3> vdd vss wl<51> / cell_PIM2
XI17192 bl<3> cbl<1> in1<50> in2<50> sl<3> vdd vss wl<50> / cell_PIM2
XI17191 bl<3> cbl<1> in1<49> in2<49> sl<3> vdd vss wl<49> / cell_PIM2
XI17190 bl<3> cbl<1> in1<48> in2<48> sl<3> vdd vss wl<48> / cell_PIM2
XI17843 bl<11> cbl<5> in1<123> in2<123> sl<11> vdd vss wl<123> / cell_PIM2
XI17842 bl<11> cbl<5> in1<124> in2<124> sl<11> vdd vss wl<124> / cell_PIM2
XI18493 bl<11> cbl<5> in1<40> in2<40> sl<11> vdd vss wl<40> / cell_PIM2
XI18492 bl<11> cbl<5> in1<41> in2<41> sl<11> vdd vss wl<41> / cell_PIM2
XI18491 bl<11> cbl<5> in1<42> in2<42> sl<11> vdd vss wl<42> / cell_PIM2
XI18490 bl<11> cbl<5> in1<43> in2<43> sl<11> vdd vss wl<43> / cell_PIM2
XI19142 bl<31> cbl<15> in1<112> in2<112> sl<31> vdd vss wl<112> / cell_PIM2
XI19143 bl<31> cbl<15> in1<111> in2<111> sl<31> vdd vss wl<111> / cell_PIM2
XI20312 bl<21> cbl<10> in1<33> in2<33> sl<21> vdd vss wl<33> / cell_PIM2
XI20311 bl<21> cbl<10> in1<32> in2<32> sl<21> vdd vss wl<32> / cell_PIM2
XI20310 bl<21> cbl<10> in1<36> in2<36> sl<21> vdd vss wl<36> / cell_PIM2
XI20309 bl<21> cbl<10> in1<35> in2<35> sl<21> vdd vss wl<35> / cell_PIM2
XI20963 bl<49> cbl<24> in1<126> in2<126> sl<49> vdd vss wl<126> / cell_PIM2
XI20962 bl<49> cbl<24> in1<125> in2<125> sl<49> vdd vss wl<125> / cell_PIM2
XI20961 bl<49> cbl<24> in1<124> in2<124> sl<49> vdd vss wl<124> / cell_PIM2
XI20960 bl<49> cbl<24> in1<123> in2<123> sl<49> vdd vss wl<123> / cell_PIM2
XI21610 bl<55> cbl<27> in1<104> in2<104> sl<55> vdd vss wl<104> / cell_PIM2
XI21609 bl<55> cbl<27> in1<105> in2<105> sl<55> vdd vss wl<105> / cell_PIM2
XI22262 bl<59> cbl<29> in1<84> in2<84> sl<59> vdd vss wl<84> / cell_PIM2
XI22261 bl<59> cbl<29> in1<85> in2<85> sl<59> vdd vss wl<85> / cell_PIM2
XI22260 bl<59> cbl<29> in1<86> in2<86> sl<59> vdd vss wl<86> / cell_PIM2
XI22259 bl<59> cbl<29> in1<87> in2<87> sl<59> vdd vss wl<87> / cell_PIM2
XI17184 bl<3> cbl<1> in1<57> in2<57> sl<3> vdd vss wl<57> / cell_PIM2
XI17834 bl<9> cbl<4> in1<122> in2<122> sl<9> vdd vss wl<122> / cell_PIM2
XI17835 bl<9> cbl<4> in1<123> in2<123> sl<9> vdd vss wl<123> / cell_PIM2
XI17836 bl<9> cbl<4> in1<124> in2<124> sl<9> vdd vss wl<124> / cell_PIM2
XI18484 bl<9> cbl<4> in1<43> in2<43> sl<9> vdd vss wl<43> / cell_PIM2
XI19134 bl<29> cbl<14> in1<108> in2<108> sl<29> vdd vss wl<108> / cell_PIM2
XI19135 bl<29> cbl<14> in1<109> in2<109> sl<29> vdd vss wl<109> / cell_PIM2
XI19136 bl<29> cbl<14> in1<110> in2<110> sl<29> vdd vss wl<110> / cell_PIM2
XI19781 bl<21> cbl<10> in1<69> in2<69> sl<21> vdd vss wl<69> / cell_PIM2
XI19782 bl<21> cbl<10> in1<65> in2<65> sl<21> vdd vss wl<65> / cell_PIM2
XI19783 bl<21> cbl<10> in1<66> in2<66> sl<21> vdd vss wl<66> / cell_PIM2
XI19784 bl<21> cbl<10> in1<67> in2<67> sl<21> vdd vss wl<67> / cell_PIM2
XI20308 bl<21> cbl<10> in1<34> in2<34> sl<21> vdd vss wl<34> / cell_PIM2
XI20954 bl<47> cbl<23> in1<127> in2<127> sl<47> vdd vss wl<127> / cell_PIM2
XI21607 bl<55> cbl<27> in1<107> in2<107> sl<55> vdd vss wl<107> / cell_PIM2
XI21608 bl<55> cbl<27> in1<106> in2<106> sl<55> vdd vss wl<106> / cell_PIM2
XI17183 bl<3> cbl<1> in1<56> in2<56> sl<3> vdd vss wl<56> / cell_PIM2
XI17182 bl<3> cbl<1> in1<55> in2<55> sl<3> vdd vss wl<55> / cell_PIM2
XI17181 bl<3> cbl<1> in1<54> in2<54> sl<3> vdd vss wl<54> / cell_PIM2
XI17180 bl<3> cbl<1> in1<53> in2<53> sl<3> vdd vss wl<53> / cell_PIM2
XI17833 bl<9> cbl<4> in1<121> in2<121> sl<9> vdd vss wl<121> / cell_PIM2
XI17832 bl<9> cbl<4> in1<120> in2<120> sl<9> vdd vss wl<120> / cell_PIM2
XI18483 bl<9> cbl<4> in1<42> in2<42> sl<9> vdd vss wl<42> / cell_PIM2
XI18482 bl<9> cbl<4> in1<41> in2<41> sl<9> vdd vss wl<41> / cell_PIM2
XI18481 bl<9> cbl<4> in1<40> in2<40> sl<9> vdd vss wl<40> / cell_PIM2
XI18480 bl<9> cbl<4> in1<39> in2<39> sl<9> vdd vss wl<39> / cell_PIM2
XI19132 bl<29> cbl<14> in1<111> in2<111> sl<29> vdd vss wl<111> / cell_PIM2
XI19133 bl<29> cbl<14> in1<112> in2<112> sl<29> vdd vss wl<112> / cell_PIM2
XI19780 bl<21> cbl<10> in1<68> in2<68> sl<21> vdd vss wl<68> / cell_PIM2
XI20302 bl<19> cbl<9> in1<32> in2<32> sl<19> vdd vss wl<32> / cell_PIM2
XI20301 bl<19> cbl<9> in1<33> in2<33> sl<19> vdd vss wl<33> / cell_PIM2
XI20300 bl<19> cbl<9> in1<34> in2<34> sl<19> vdd vss wl<34> / cell_PIM2
XI20299 bl<19> cbl<9> in1<35> in2<35> sl<19> vdd vss wl<35> / cell_PIM2
XI20953 bl<47> cbl<23> in1<126> in2<126> sl<47> vdd vss wl<126> / cell_PIM2
XI20952 bl<47> cbl<23> in1<125> in2<125> sl<47> vdd vss wl<125> / cell_PIM2
XI20951 bl<47> cbl<23> in1<123> in2<123> sl<47> vdd vss wl<123> / cell_PIM2
XI20950 bl<47> cbl<23> in1<124> in2<124> sl<47> vdd vss wl<124> / cell_PIM2
XI21602 bl<53> cbl<26> in1<105> in2<105> sl<53> vdd vss wl<105> / cell_PIM2
XI21601 bl<53> cbl<26> in1<104> in2<104> sl<53> vdd vss wl<104> / cell_PIM2
XI21600 bl<53> cbl<26> in1<107> in2<107> sl<53> vdd vss wl<107> / cell_PIM2
XI21599 bl<53> cbl<26> in1<106> in2<106> sl<53> vdd vss wl<106> / cell_PIM2
XI22252 bl<57> cbl<28> in1<84> in2<84> sl<57> vdd vss wl<84> / cell_PIM2
XI22251 bl<57> cbl<28> in1<85> in2<85> sl<57> vdd vss wl<85> / cell_PIM2
XI22250 bl<57> cbl<28> in1<86> in2<86> sl<57> vdd vss wl<86> / cell_PIM2
XI22249 bl<57> cbl<28> in1<87> in2<87> sl<57> vdd vss wl<87> / cell_PIM2
XI22898 bl<33> cbl<16> in1<62> in2<62> sl<33> vdd vss wl<62> / cell_PIM2
XI22897 bl<33> cbl<16> in1<61> in2<61> sl<33> vdd vss wl<61> / cell_PIM2
XI24072 bl<57> cbl<28> in1<31> in2<31> sl<57> vdd vss wl<31> / cell_PIM2
XI24073 bl<57> cbl<28> in1<30> in2<30> sl<57> vdd vss wl<30> / cell_PIM2
XI24722 bl<33> cbl<16> in1<7> in2<7> sl<33> vdd vss wl<7> / cell_PIM2
XI24721 bl<33> cbl<16> in1<6> in2<6> sl<33> vdd vss wl<6> / cell_PIM2
XI24720 bl<33> cbl<16> in1<5> in2<5> sl<33> vdd vss wl<5> / cell_PIM2
XI24723 bl<33> cbl<16> in1<4> in2<4> sl<33> vdd vss wl<4> / cell_PIM2
XI17174 bl<3> cbl<1> in1<62> in2<62> sl<3> vdd vss wl<62> / cell_PIM2
XI17826 bl<15> cbl<7> in1<127> in2<127> sl<15> vdd vss wl<127> / cell_PIM2
XI17825 bl<15> cbl<7> in1<126> in2<126> sl<15> vdd vss wl<126> / cell_PIM2
XI17824 bl<15> cbl<7> in1<125> in2<125> sl<15> vdd vss wl<125> / cell_PIM2
XI18474 bl<15> cbl<7> in1<44> in2<44> sl<15> vdd vss wl<44> / cell_PIM2
XI19126 bl<27> cbl<13> in1<108> in2<108> sl<27> vdd vss wl<108> / cell_PIM2
XI19125 bl<27> cbl<13> in1<109> in2<109> sl<27> vdd vss wl<109> / cell_PIM2
XI19124 bl<27> cbl<13> in1<110> in2<110> sl<27> vdd vss wl<110> / cell_PIM2
XI19774 bl<19> cbl<9> in1<65> in2<65> sl<19> vdd vss wl<65> / cell_PIM2
XI19773 bl<19> cbl<9> in1<66> in2<66> sl<19> vdd vss wl<66> / cell_PIM2
XI20298 bl<19> cbl<9> in1<36> in2<36> sl<19> vdd vss wl<36> / cell_PIM2
XI20944 bl<45> cbl<22> in1<127> in2<127> sl<45> vdd vss wl<127> / cell_PIM2
XI21594 bl<51> cbl<25> in1<104> in2<104> sl<51> vdd vss wl<104> / cell_PIM2
XI22248 bl<57> cbl<28> in1<88> in2<88> sl<57> vdd vss wl<88> / cell_PIM2
XI22896 bl<33> cbl<16> in1<64> in2<64> sl<33> vdd vss wl<64> / cell_PIM2
XI22895 bl<33> cbl<16> in1<63> in2<63> sl<33> vdd vss wl<63> / cell_PIM2
XI23418 bl<47> cbl<23> in1<46> in2<46> sl<47> vdd vss wl<46> / cell_PIM2
XI23417 bl<47> cbl<23> in1<47> in2<47> sl<47> vdd vss wl<47> / cell_PIM2
XI23416 bl<47> cbl<23> in1<48> in2<48> sl<47> vdd vss wl<48> / cell_PIM2
XI23415 bl<47> cbl<23> in1<49> in2<49> sl<47> vdd vss wl<49> / cell_PIM2
XI23414 bl<47> cbl<23> in1<50> in2<50> sl<47> vdd vss wl<50> / cell_PIM2
XI24066 bl<55> cbl<27> in1<27> in2<27> sl<55> vdd vss wl<27> / cell_PIM2
XI24065 bl<55> cbl<27> in1<28> in2<28> sl<55> vdd vss wl<28> / cell_PIM2
XI24064 bl<55> cbl<27> in1<29> in2<29> sl<55> vdd vss wl<29> / cell_PIM2
XI24714 bl<63> cbl<31> in1<8> in2<8> sl<63> vdd vss wl<8> / cell_PIM2
XI16908 bl<1> cbl<0> in1<1> in2<1> sl<1> vdd vss wl<1> / cell_PIM2
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv8
* View Name:    schematic
************************************************************************

.SUBCKT inv8 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=1u
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=1u
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    nand
* View Name:    schematic
************************************************************************

.SUBCKT nand IN0 IN1 OUT VDD VSS
*.PININFO IN0:B IN1:B OUT:B VDD:B VSS:B
XNM4 net10 IN1 VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM3 OUT IN0 net10 VSS n12ll_mis_ckt MR=1 L=60n W=120n
XPM2 OUT IN1 VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM1 OUT IN0 VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    mux8x1
* View Name:    schematic
************************************************************************

.SUBCKT mux8x1 group<0> group<1> group<2> group<3> group<4> group<5> group<6> 
+ group<7> in out<0> out<1> out<2> out<3> out<4> out<5> out<6> out<7> vdd vss
*.PININFO group<0>:I group<1>:I group<2>:I group<3>:I group<4>:I group<5>:I 
*.PININFO group<6>:I group<7>:I in:I out<0>:O out<1>:O out<2>:O out<3>:O 
*.PININFO out<4>:O out<5>:O out<6>:O out<7>:O vdd:B vss:B
XI19 net80 out<0> vdd vss / inv8
XI17 net81 out<1> vdd vss / inv8
XI6 net82 out<2> vdd vss / inv8
XI7 net83 out<3> vdd vss / inv8
XI9 net84 out<4> vdd vss / inv8
XI11 net85 out<5> vdd vss / inv8
XI13 net86 out<6> vdd vss / inv8
XI15 net87 out<7> vdd vss / inv8
XI23 in group<0> net80 vdd vss / nand
XI22 in group<1> net81 vdd vss / nand
XI21 in group<2> net82 vdd vss / nand
XI4 in group<7> net87 vdd vss / nand
XI0 in group<3> net83 vdd vss / nand
XI1 in group<4> net84 vdd vss / nand
XI2 in group<5> net85 vdd vss / nand
XI3 in group<6> net86 vdd vss / nand
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    WLdriver
* View Name:    schematic
************************************************************************

.SUBCKT WLdriver blbuf<0> blbuf<1> blbuf<2> blbuf<3> blbuf<4> blbuf<5> 
+ blbuf<6> blbuf<7> blbuf<8> blbuf<9> blbuf<10> blbuf<11> blbuf<12> blbuf<13> 
+ blbuf<14> blbuf<15> group<0> group<1> group<2> group<3> group<4> group<5> 
+ group<6> group<7> in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> in1<7> 
+ in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> 
+ in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> 
+ in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> 
+ in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> 
+ in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> 
+ in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> 
+ in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> 
+ in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> 
+ in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> 
+ in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> 
+ in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> 
+ in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> in1<113> 
+ in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> 
+ in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> in2<2> 
+ in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> 
+ in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> 
+ in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> 
+ in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> in2<39> 
+ in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> in2<48> 
+ in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> in2<57> 
+ in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> in2<66> 
+ in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> 
+ in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> in2<84> 
+ in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> 
+ in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> in2<102> 
+ in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> in2<110> 
+ in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> in2<118> 
+ in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> in2<126> 
+ in2<127> row16<0> row16<1> row16<2> row16<3> row16<4> row16<5> row16<6> 
+ row16<7> row16<8> row16<9> row16<10> row16<11> row16<12> row16<13> row16<14> 
+ row16<15> slbuf<0> slbuf<1> slbuf<2> slbuf<3> slbuf<4> slbuf<5> slbuf<6> 
+ slbuf<7> slbuf<8> slbuf<9> slbuf<10> slbuf<11> slbuf<12> slbuf<13> slbuf<14> 
+ slbuf<15> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> 
+ wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> 
+ wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> 
+ wl<31> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> wl<40> wl<41> 
+ wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> wl<48> wl<49> wl<50> wl<51> wl<52> 
+ wl<53> wl<54> wl<55> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> 
+ wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> wl<72> wl<73> wl<74> 
+ wl<75> wl<76> wl<77> wl<78> wl<79> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> 
+ wl<86> wl<87> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> wl<96> 
+ wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> wl<104> wl<105> wl<106> 
+ wl<107> wl<108> wl<109> wl<110> wl<111> wl<112> wl<113> wl<114> wl<115> 
+ wl<116> wl<117> wl<118> wl<119> wl<120> wl<121> wl<122> wl<123> wl<124> 
+ wl<125> wl<126> wl<127>
*.PININFO group<0>:I group<1>:I group<2>:I group<3>:I group<4>:I group<5>:I 
*.PININFO group<6>:I group<7>:I row16<0>:I row16<1>:I row16<2>:I row16<3>:I 
*.PININFO row16<4>:I row16<5>:I row16<6>:I row16<7>:I row16<8>:I row16<9>:I 
*.PININFO row16<10>:I row16<11>:I row16<12>:I row16<13>:I row16<14>:I 
*.PININFO row16<15>:I wl<0>:O wl<1>:O wl<2>:O wl<3>:O wl<4>:O wl<5>:O wl<6>:O 
*.PININFO wl<7>:O wl<8>:O wl<9>:O wl<10>:O wl<11>:O wl<12>:O wl<13>:O wl<14>:O 
*.PININFO wl<15>:O wl<16>:O wl<17>:O wl<18>:O wl<19>:O wl<20>:O wl<21>:O 
*.PININFO wl<22>:O wl<23>:O wl<24>:O wl<25>:O wl<26>:O wl<27>:O wl<28>:O 
*.PININFO wl<29>:O wl<30>:O wl<31>:O wl<32>:O wl<33>:O wl<34>:O wl<35>:O 
*.PININFO wl<36>:O wl<37>:O wl<38>:O wl<39>:O wl<40>:O wl<41>:O wl<42>:O 
*.PININFO wl<43>:O wl<44>:O wl<45>:O wl<46>:O wl<47>:O wl<48>:O wl<49>:O 
*.PININFO wl<50>:O wl<51>:O wl<52>:O wl<53>:O wl<54>:O wl<55>:O wl<56>:O 
*.PININFO wl<57>:O wl<58>:O wl<59>:O wl<60>:O wl<61>:O wl<62>:O wl<63>:O 
*.PININFO wl<64>:O wl<65>:O wl<66>:O wl<67>:O wl<68>:O wl<69>:O wl<70>:O 
*.PININFO wl<71>:O wl<72>:O wl<73>:O wl<74>:O wl<75>:O wl<76>:O wl<77>:O 
*.PININFO wl<78>:O wl<79>:O wl<80>:O wl<81>:O wl<82>:O wl<83>:O wl<84>:O 
*.PININFO wl<85>:O wl<86>:O wl<87>:O wl<88>:O wl<89>:O wl<90>:O wl<91>:O 
*.PININFO wl<92>:O wl<93>:O wl<94>:O wl<95>:O wl<96>:O wl<97>:O wl<98>:O 
*.PININFO wl<99>:O wl<100>:O wl<101>:O wl<102>:O wl<103>:O wl<104>:O wl<105>:O 
*.PININFO wl<106>:O wl<107>:O wl<108>:O wl<109>:O wl<110>:O wl<111>:O 
*.PININFO wl<112>:O wl<113>:O wl<114>:O wl<115>:O wl<116>:O wl<117>:O 
*.PININFO wl<118>:O wl<119>:O wl<120>:O wl<121>:O wl<122>:O wl<123>:O 
*.PININFO wl<124>:O wl<125>:O wl<126>:O wl<127>:O blbuf<0>:B blbuf<1>:B 
*.PININFO blbuf<2>:B blbuf<3>:B blbuf<4>:B blbuf<5>:B blbuf<6>:B blbuf<7>:B 
*.PININFO blbuf<8>:B blbuf<9>:B blbuf<10>:B blbuf<11>:B blbuf<12>:B 
*.PININFO blbuf<13>:B blbuf<14>:B blbuf<15>:B in1<0>:B in1<1>:B in1<2>:B 
*.PININFO in1<3>:B in1<4>:B in1<5>:B in1<6>:B in1<7>:B in1<8>:B in1<9>:B 
*.PININFO in1<10>:B in1<11>:B in1<12>:B in1<13>:B in1<14>:B in1<15>:B 
*.PININFO in1<16>:B in1<17>:B in1<18>:B in1<19>:B in1<20>:B in1<21>:B 
*.PININFO in1<22>:B in1<23>:B in1<24>:B in1<25>:B in1<26>:B in1<27>:B 
*.PININFO in1<28>:B in1<29>:B in1<30>:B in1<31>:B in1<32>:B in1<33>:B 
*.PININFO in1<34>:B in1<35>:B in1<36>:B in1<37>:B in1<38>:B in1<39>:B 
*.PININFO in1<40>:B in1<41>:B in1<42>:B in1<43>:B in1<44>:B in1<45>:B 
*.PININFO in1<46>:B in1<47>:B in1<48>:B in1<49>:B in1<50>:B in1<51>:B 
*.PININFO in1<52>:B in1<53>:B in1<54>:B in1<55>:B in1<56>:B in1<57>:B 
*.PININFO in1<58>:B in1<59>:B in1<60>:B in1<61>:B in1<62>:B in1<63>:B 
*.PININFO in1<64>:B in1<65>:B in1<66>:B in1<67>:B in1<68>:B in1<69>:B 
*.PININFO in1<70>:B in1<71>:B in1<72>:B in1<73>:B in1<74>:B in1<75>:B 
*.PININFO in1<76>:B in1<77>:B in1<78>:B in1<79>:B in1<80>:B in1<81>:B 
*.PININFO in1<82>:B in1<83>:B in1<84>:B in1<85>:B in1<86>:B in1<87>:B 
*.PININFO in1<88>:B in1<89>:B in1<90>:B in1<91>:B in1<92>:B in1<93>:B 
*.PININFO in1<94>:B in1<95>:B in1<96>:B in1<97>:B in1<98>:B in1<99>:B 
*.PININFO in1<100>:B in1<101>:B in1<102>:B in1<103>:B in1<104>:B in1<105>:B 
*.PININFO in1<106>:B in1<107>:B in1<108>:B in1<109>:B in1<110>:B in1<111>:B 
*.PININFO in1<112>:B in1<113>:B in1<114>:B in1<115>:B in1<116>:B in1<117>:B 
*.PININFO in1<118>:B in1<119>:B in1<120>:B in1<121>:B in1<122>:B in1<123>:B 
*.PININFO in1<124>:B in1<125>:B in1<126>:B in1<127>:B in2<0>:B in2<1>:B 
*.PININFO in2<2>:B in2<3>:B in2<4>:B in2<5>:B in2<6>:B in2<7>:B in2<8>:B 
*.PININFO in2<9>:B in2<10>:B in2<11>:B in2<12>:B in2<13>:B in2<14>:B in2<15>:B 
*.PININFO in2<16>:B in2<17>:B in2<18>:B in2<19>:B in2<20>:B in2<21>:B 
*.PININFO in2<22>:B in2<23>:B in2<24>:B in2<25>:B in2<26>:B in2<27>:B 
*.PININFO in2<28>:B in2<29>:B in2<30>:B in2<31>:B in2<32>:B in2<33>:B 
*.PININFO in2<34>:B in2<35>:B in2<36>:B in2<37>:B in2<38>:B in2<39>:B 
*.PININFO in2<40>:B in2<41>:B in2<42>:B in2<43>:B in2<44>:B in2<45>:B 
*.PININFO in2<46>:B in2<47>:B in2<48>:B in2<49>:B in2<50>:B in2<51>:B 
*.PININFO in2<52>:B in2<53>:B in2<54>:B in2<55>:B in2<56>:B in2<57>:B 
*.PININFO in2<58>:B in2<59>:B in2<60>:B in2<61>:B in2<62>:B in2<63>:B 
*.PININFO in2<64>:B in2<65>:B in2<66>:B in2<67>:B in2<68>:B in2<69>:B 
*.PININFO in2<70>:B in2<71>:B in2<72>:B in2<73>:B in2<74>:B in2<75>:B 
*.PININFO in2<76>:B in2<77>:B in2<78>:B in2<79>:B in2<80>:B in2<81>:B 
*.PININFO in2<82>:B in2<83>:B in2<84>:B in2<85>:B in2<86>:B in2<87>:B 
*.PININFO in2<88>:B in2<89>:B in2<90>:B in2<91>:B in2<92>:B in2<93>:B 
*.PININFO in2<94>:B in2<95>:B in2<96>:B in2<97>:B in2<98>:B in2<99>:B 
*.PININFO in2<100>:B in2<101>:B in2<102>:B in2<103>:B in2<104>:B in2<105>:B 
*.PININFO in2<106>:B in2<107>:B in2<108>:B in2<109>:B in2<110>:B in2<111>:B 
*.PININFO in2<112>:B in2<113>:B in2<114>:B in2<115>:B in2<116>:B in2<117>:B 
*.PININFO in2<118>:B in2<119>:B in2<120>:B in2<121>:B in2<122>:B in2<123>:B 
*.PININFO in2<124>:B in2<125>:B in2<126>:B in2<127>:B slbuf<0>:B slbuf<1>:B 
*.PININFO slbuf<2>:B slbuf<3>:B slbuf<4>:B slbuf<5>:B slbuf<6>:B slbuf<7>:B 
*.PININFO slbuf<8>:B slbuf<9>:B slbuf<10>:B slbuf<11>:B slbuf<12>:B 
*.PININFO slbuf<13>:B slbuf<14>:B slbuf<15>:B vdd:B vss:B
XI16 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<15> wl<120> wl<121> wl<122> wl<123> wl<124> wl<125> wl<126> wl<127> 
+ vdd vss / mux8x1
XI15 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<14> wl<112> wl<113> wl<114> wl<115> wl<116> wl<117> wl<118> wl<119> 
+ vdd vss / mux8x1
XI14 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<13> wl<104> wl<105> wl<106> wl<107> wl<108> wl<109> wl<110> wl<111> 
+ vdd vss / mux8x1
XI13 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<12> wl<96> wl<97> wl<98> wl<99> wl<100> wl<101> wl<102> wl<103> vdd 
+ vss / mux8x1
XI12 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<11> wl<88> wl<89> wl<90> wl<91> wl<92> wl<93> wl<94> wl<95> vdd vss / 
+ mux8x1
XI11 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<10> wl<80> wl<81> wl<82> wl<83> wl<84> wl<85> wl<86> wl<87> vdd vss / 
+ mux8x1
XI10 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<9> wl<72> wl<73> wl<74> wl<75> wl<76> wl<77> wl<78> wl<79> vdd vss / 
+ mux8x1
XI9 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<8> wl<64> wl<65> wl<66> wl<67> wl<68> wl<69> wl<70> wl<71> vdd vss / 
+ mux8x1
XI8 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<7> wl<56> wl<57> wl<58> wl<59> wl<60> wl<61> wl<62> wl<63> vdd vss / 
+ mux8x1
XI7 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<6> wl<48> wl<49> wl<50> wl<51> wl<52> wl<53> wl<54> wl<55> vdd vss / 
+ mux8x1
XI6 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<5> wl<40> wl<41> wl<42> wl<43> wl<44> wl<45> wl<46> wl<47> vdd vss / 
+ mux8x1
XI5 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<4> wl<32> wl<33> wl<34> wl<35> wl<36> wl<37> wl<38> wl<39> vdd vss / 
+ mux8x1
XI4 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<3> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> vdd vss / 
+ mux8x1
XI1 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<0> wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> vdd vss / mux8x1
XI2 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<1> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> vdd vss / 
+ mux8x1
XI3 group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<2> wl<16> wl<17> wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> vdd vss / 
+ mux8x1
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    nor
* View Name:    schematic
************************************************************************

.SUBCKT nor IN0 IN1 OUT VDD VSS
*.PININFO IN0:B IN1:B OUT:B VDD:B VSS:B
XNM2 OUT IN1 VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM3 OUT IN0 VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XPM3 OUT IN1 net018 VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM0 net018 IN0 VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv2
* View Name:    schematic
************************************************************************

.SUBCKT inv2 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=60n W=900n
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=60n W=1.8u
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    Tgate
* View Name:    schematic
************************************************************************

.SUBCKT Tgate IN OE OEN OUT VDD VSS
*.PININFO IN:B OE:B OEN:B OUT:B VDD:B VSS:B
XNM2 OUT OE IN VSS n12ll_mis_ckt MR=1 L=60n W=600n
XPM0 IN OEN OUT VDD p12ll_mis_ckt MR=1 L=60n W=1.2u
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv1
* View Name:    schematic
************************************************************************

.SUBCKT inv1 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=60n W=900n
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=60n W=450n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Writecell
* View Name:    schematic
************************************************************************

.SUBCKT Writecell VDD VSS bl<0> bl<1> bl<2> bl<3> blbuf col<0> col<1> col<2> 
+ col<3> d sl<0> sl<1> sl<2> sl<3> slbuf wrt wrtbuf
*.PININFO col<0>:I col<1>:I col<2>:I col<3>:I d:I wrt:I wrtbuf:I bl<0>:O 
*.PININFO bl<1>:O bl<2>:O bl<3>:O blbuf:O sl<0>:O sl<1>:O sl<2>:O sl<3>:O 
*.PININFO slbuf:O VDD:B VSS:B
XI15 wrt wrtbuf net013 VDD VSS / nor
XI12 wrtalln d wdnb VDD VSS / nor
XI5 wrtalln dn wdns VDD VSS / nor
XI13 wdnb wdps VDD VSS / inv2
XI6 wdns wdpb VDD VSS / inv2
XI7 d dn VDD VSS / inv2
XI3<0> wrt col<0> net042<0> VDD VSS / nand
XI3<1> wrt col<1> net042<1> VDD VSS / nand
XI3<2> wrt col<2> net042<2> VDD VSS / nand
XI3<3> wrt col<3> net042<3> VDD VSS / nand
XI19 blbuf net012 net015 tBL VDD VSS / Tgate
XI20 slbuf net012 net015 tSL VDD VSS / Tgate
XI10<0> sl<0> net043<0> net044<0> tSL VDD VSS / Tgate
XI10<1> sl<1> net043<1> net044<1> tSL VDD VSS / Tgate
XI10<2> sl<2> net043<2> net044<2> tSL VDD VSS / Tgate
XI10<3> sl<3> net043<3> net044<3> tSL VDD VSS / Tgate
XI9<0> bl<0> net043<0> net044<0> tBL VDD VSS / Tgate
XI9<1> bl<1> net043<1> net044<1> tBL VDD VSS / Tgate
XI9<2> bl<2> net043<2> net044<2> tBL VDD VSS / Tgate
XI9<3> bl<3> net043<3> net044<3> tBL VDD VSS / Tgate
XI22 wrtbuf net024 VDD VSS / inv1
XI17 net024 net012 VDD VSS / inv1
XI21 net012 net015 VDD VSS / inv1
XI16 net013 wrtall VDD VSS / inv1
XI8<0> net043<0> net044<0> VDD VSS / inv1
XI8<1> net043<1> net044<1> VDD VSS / inv1
XI8<2> net043<2> net044<2> VDD VSS / inv1
XI8<3> net043<3> net044<3> VDD VSS / inv1
XI11 wrtall wrtalln VDD VSS / inv1
XI14<0> net042<0> net043<0> VDD VSS / inv1
XI14<1> net042<1> net043<1> VDD VSS / inv1
XI14<2> net042<2> net043<2> VDD VSS / inv1
XI14<3> net042<3> net043<3> VDD VSS / inv1
XPM2 tBL wdpb VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XPM1 tSL wdps VDD VDD p12ll_mis_ckt MR=1 L=60n W=120n
XNM0 tBL wdnb VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
XNM1 tSL wdns VSS VSS n12ll_mis_ckt MR=1 L=60n W=120n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Writedriver
* View Name:    schematic
************************************************************************

.SUBCKT Writedriver bl<0> bl<1> bl<2> bl<3> bl<4> bl<5> bl<6> bl<7> bl<8> 
+ bl<9> bl<10> bl<11> bl<12> bl<13> bl<14> bl<15> bl<16> bl<17> bl<18> bl<19> 
+ bl<20> bl<21> bl<22> bl<23> bl<24> bl<25> bl<26> bl<27> bl<28> bl<29> bl<30> 
+ bl<31> bl<32> bl<33> bl<34> bl<35> bl<36> bl<37> bl<38> bl<39> bl<40> bl<41> 
+ bl<42> bl<43> bl<44> bl<45> bl<46> bl<47> bl<48> bl<49> bl<50> bl<51> bl<52> 
+ bl<53> bl<54> bl<55> bl<56> bl<57> bl<58> bl<59> bl<60> bl<61> bl<62> bl<63> 
+ blbuf<0> blbuf<1> blbuf<2> blbuf<3> blbuf<4> blbuf<5> blbuf<6> blbuf<7> 
+ blbuf<8> blbuf<9> blbuf<10> blbuf<11> blbuf<12> blbuf<13> blbuf<14> 
+ blbuf<15> cbl<0> cbl<1> cbl<2> cbl<3> cbl<4> cbl<5> cbl<6> cbl<7> cbl<8> 
+ cbl<9> cbl<10> cbl<11> cbl<12> cbl<13> cbl<14> cbl<15> cbl<16> cbl<17> 
+ cbl<18> cbl<19> cbl<20> cbl<21> cbl<22> cbl<23> cbl<24> cbl<25> cbl<26> 
+ cbl<27> cbl<28> cbl<29> cbl<30> cbl<31> col<0> col<1> col<2> col<3> d<0> 
+ d<1> d<2> d<3> d<4> d<5> d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> 
+ d<15> sl<0> sl<1> sl<2> sl<3> sl<4> sl<5> sl<6> sl<7> sl<8> sl<9> sl<10> 
+ sl<11> sl<12> sl<13> sl<14> sl<15> sl<16> sl<17> sl<18> sl<19> sl<20> sl<21> 
+ sl<22> sl<23> sl<24> sl<25> sl<26> sl<27> sl<28> sl<29> sl<30> sl<31> sl<32> 
+ sl<33> sl<34> sl<35> sl<36> sl<37> sl<38> sl<39> sl<40> sl<41> sl<42> sl<43> 
+ sl<44> sl<45> sl<46> sl<47> sl<48> sl<49> sl<50> sl<51> sl<52> sl<53> sl<54> 
+ sl<55> sl<56> sl<57> sl<58> sl<59> sl<60> sl<61> sl<62> sl<63> slbuf<0> 
+ slbuf<1> slbuf<2> slbuf<3> slbuf<4> slbuf<5> slbuf<6> slbuf<7> slbuf<8> 
+ slbuf<9> slbuf<10> slbuf<11> slbuf<12> slbuf<13> slbuf<14> slbuf<15> vdd vss 
+ wrt wrtbuf
*.PININFO col<0>:I col<1>:I col<2>:I col<3>:I d<0>:I d<1>:I d<2>:I d<3>:I 
*.PININFO d<4>:I d<5>:I d<6>:I d<7>:I d<8>:I d<9>:I d<10>:I d<11>:I d<12>:I 
*.PININFO d<13>:I d<14>:I d<15>:I wrt:I wrtbuf:I bl<0>:O bl<1>:O bl<2>:O 
*.PININFO bl<3>:O bl<4>:O bl<5>:O bl<6>:O bl<7>:O bl<8>:O bl<9>:O bl<10>:O 
*.PININFO bl<11>:O bl<12>:O bl<13>:O bl<14>:O bl<15>:O bl<16>:O bl<17>:O 
*.PININFO bl<18>:O bl<19>:O bl<20>:O bl<21>:O bl<22>:O bl<23>:O bl<24>:O 
*.PININFO bl<25>:O bl<26>:O bl<27>:O bl<28>:O bl<29>:O bl<30>:O bl<31>:O 
*.PININFO bl<32>:O bl<33>:O bl<34>:O bl<35>:O bl<36>:O bl<37>:O bl<38>:O 
*.PININFO bl<39>:O bl<40>:O bl<41>:O bl<42>:O bl<43>:O bl<44>:O bl<45>:O 
*.PININFO bl<46>:O bl<47>:O bl<48>:O bl<49>:O bl<50>:O bl<51>:O bl<52>:O 
*.PININFO bl<53>:O bl<54>:O bl<55>:O bl<56>:O bl<57>:O bl<58>:O bl<59>:O 
*.PININFO bl<60>:O bl<61>:O bl<62>:O bl<63>:O blbuf<0>:O blbuf<1>:O blbuf<2>:O 
*.PININFO blbuf<3>:O blbuf<4>:O blbuf<5>:O blbuf<6>:O blbuf<7>:O blbuf<8>:O 
*.PININFO blbuf<9>:O blbuf<10>:O blbuf<11>:O blbuf<12>:O blbuf<13>:O 
*.PININFO blbuf<14>:O blbuf<15>:O sl<0>:O sl<1>:O sl<2>:O sl<3>:O sl<4>:O 
*.PININFO sl<5>:O sl<6>:O sl<7>:O sl<8>:O sl<9>:O sl<10>:O sl<11>:O sl<12>:O 
*.PININFO sl<13>:O sl<14>:O sl<15>:O sl<16>:O sl<17>:O sl<18>:O sl<19>:O 
*.PININFO sl<20>:O sl<21>:O sl<22>:O sl<23>:O sl<24>:O sl<25>:O sl<26>:O 
*.PININFO sl<27>:O sl<28>:O sl<29>:O sl<30>:O sl<31>:O sl<32>:O sl<33>:O 
*.PININFO sl<34>:O sl<35>:O sl<36>:O sl<37>:O sl<38>:O sl<39>:O sl<40>:O 
*.PININFO sl<41>:O sl<42>:O sl<43>:O sl<44>:O sl<45>:O sl<46>:O sl<47>:O 
*.PININFO sl<48>:O sl<49>:O sl<50>:O sl<51>:O sl<52>:O sl<53>:O sl<54>:O 
*.PININFO sl<55>:O sl<56>:O sl<57>:O sl<58>:O sl<59>:O sl<60>:O sl<61>:O 
*.PININFO sl<62>:O sl<63>:O slbuf<0>:O slbuf<1>:O slbuf<2>:O slbuf<3>:O 
*.PININFO slbuf<4>:O slbuf<5>:O slbuf<6>:O slbuf<7>:O slbuf<8>:O slbuf<9>:O 
*.PININFO slbuf<10>:O slbuf<11>:O slbuf<12>:O slbuf<13>:O slbuf<14>:O 
*.PININFO slbuf<15>:O cbl<0>:B cbl<1>:B cbl<2>:B cbl<3>:B cbl<4>:B cbl<5>:B 
*.PININFO cbl<6>:B cbl<7>:B cbl<8>:B cbl<9>:B cbl<10>:B cbl<11>:B cbl<12>:B 
*.PININFO cbl<13>:B cbl<14>:B cbl<15>:B cbl<16>:B cbl<17>:B cbl<18>:B 
*.PININFO cbl<19>:B cbl<20>:B cbl<21>:B cbl<22>:B cbl<23>:B cbl<24>:B 
*.PININFO cbl<25>:B cbl<26>:B cbl<27>:B cbl<28>:B cbl<29>:B cbl<30>:B 
*.PININFO cbl<31>:B vdd:B vss:B
XI16 vdd vss bl<60> bl<61> bl<62> bl<63> blbuf<15> col<0> col<1> col<2> col<3> 
+ d<15> sl<60> sl<61> sl<62> sl<63> slbuf<15> wrt wrtbuf / Writecell
XI15 vdd vss bl<56> bl<57> bl<58> bl<59> blbuf<14> col<0> col<1> col<2> col<3> 
+ d<14> sl<56> sl<57> sl<58> sl<59> slbuf<14> wrt wrtbuf / Writecell
XI14 vdd vss bl<52> bl<53> bl<54> bl<55> blbuf<13> col<0> col<1> col<2> col<3> 
+ d<13> sl<52> sl<53> sl<54> sl<55> slbuf<13> wrt wrtbuf / Writecell
XI13 vdd vss bl<48> bl<49> bl<50> bl<51> blbuf<12> col<0> col<1> col<2> col<3> 
+ d<12> sl<48> sl<49> sl<50> sl<51> slbuf<12> wrt wrtbuf / Writecell
XI12 vdd vss bl<44> bl<45> bl<46> bl<47> blbuf<11> col<0> col<1> col<2> col<3> 
+ d<11> sl<44> sl<45> sl<46> sl<47> slbuf<11> wrt wrtbuf / Writecell
XI11 vdd vss bl<40> bl<41> bl<42> bl<43> blbuf<10> col<0> col<1> col<2> col<3> 
+ d<10> sl<40> sl<41> sl<42> sl<43> slbuf<10> wrt wrtbuf / Writecell
XI10 vdd vss bl<36> bl<37> bl<38> bl<39> blbuf<9> col<0> col<1> col<2> col<3> 
+ d<9> sl<36> sl<37> sl<38> sl<39> slbuf<9> wrt wrtbuf / Writecell
XI9 vdd vss bl<32> bl<33> bl<34> bl<35> blbuf<8> col<0> col<1> col<2> col<3> 
+ d<8> sl<32> sl<33> sl<34> sl<35> slbuf<8> wrt wrtbuf / Writecell
XI8 vdd vss bl<28> bl<29> bl<30> bl<31> blbuf<7> col<0> col<1> col<2> col<3> 
+ d<7> sl<28> sl<29> sl<30> sl<31> slbuf<7> wrt wrtbuf / Writecell
XI7 vdd vss bl<24> bl<25> bl<26> bl<27> blbuf<6> col<0> col<1> col<2> col<3> 
+ d<6> sl<24> sl<25> sl<26> sl<27> slbuf<6> wrt wrtbuf / Writecell
XI6 vdd vss bl<20> bl<21> bl<22> bl<23> blbuf<5> col<0> col<1> col<2> col<3> 
+ d<5> sl<20> sl<21> sl<22> sl<23> slbuf<5> wrt wrtbuf / Writecell
XI5 vdd vss bl<16> bl<17> bl<18> bl<19> blbuf<4> col<0> col<1> col<2> col<3> 
+ d<4> sl<16> sl<17> sl<18> sl<19> slbuf<4> wrt wrtbuf / Writecell
XI4 vdd vss bl<12> bl<13> bl<14> bl<15> blbuf<3> col<0> col<1> col<2> col<3> 
+ d<3> sl<12> sl<13> sl<14> sl<15> slbuf<3> wrt wrtbuf / Writecell
XI3 vdd vss bl<8> bl<9> bl<10> bl<11> blbuf<2> col<0> col<1> col<2> col<3> 
+ d<2> sl<8> sl<9> sl<10> sl<11> slbuf<2> wrt wrtbuf / Writecell
XI2 vdd vss bl<4> bl<5> bl<6> bl<7> blbuf<1> col<0> col<1> col<2> col<3> d<1> 
+ sl<4> sl<5> sl<6> sl<7> slbuf<1> wrt wrtbuf / Writecell
XI1 vdd vss bl<0> bl<1> bl<2> bl<3> blbuf<0> col<0> col<1> col<2> col<3> d<0> 
+ sl<0> sl<1> sl<2> sl<3> slbuf<0> wrt wrtbuf / Writecell
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    3nand
* View Name:    schematic
************************************************************************

.SUBCKT 3nand VDD VSS in<0> in<1> in<2> out
*.PININFO in<0>:I in<1>:I in<2>:I out:O VDD:B VSS:B
XPM0 out in<0> VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XPM1 out in<2> VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XPM2 out in<1> VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XNM6 net12 in<2> VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
XNM5 net19 in<1> net12 VSS n12ll_mis_ckt MR=1 L=80n W=200n
XNM4 out in<0> net19 VSS n12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv4
* View Name:    schematic
************************************************************************

.SUBCKT inv4 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=60n W=1.8u
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=60n W=3.6u
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    2x4decoder
* View Name:    schematic
************************************************************************

.SUBCKT 2x4decoder VDD VSS en in<0> in<1> nout<0> nout<1> nout<2> nout<3>
*.PININFO en:I in<0>:I in<1>:I nout<0>:O nout<1>:O nout<2>:O nout<3>:O VDD:B 
*.PININFO VSS:B
XI3 VDD VSS in<0> net06 in<1> net016 / 3nand
XI2 VDD VSS net11 net06 in<1> net017 / 3nand
XI1 VDD VSS in<0> net06 net04 net018 / 3nand
XI0 VDD VSS net11 net06 net04 net019 / 3nand
XI6 en net06 VDD VSS / inv1
XI5 in<1> net04 VDD VSS / inv1
XI4 in<0> net11 VDD VSS / inv1
XI44 net016 nout<3> VDD VSS / inv4
XI43 net017 nout<2> VDD VSS / inv4
XI42 net018 nout<1> VDD VSS / inv4
XI41 net019 nout<0> VDD VSS / inv4
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    3x8decoder
* View Name:    schematic
************************************************************************

.SUBCKT 3x8decoder in<0> in<1> in<2> out<0> out<1> out<2> out<3> out<4> out<5> 
+ out<6> out<7> vdd vss
*.PININFO in<0>:I in<1>:I in<2>:I out<0>:O out<1>:O out<2>:O out<3>:O out<4>:O 
*.PININFO out<5>:O out<6>:O out<7>:O vdd:B vss:B
XI1 vdd vss inn<2> in<0> in<1> out<4> out<5> out<6> out<7> / 2x4decoder
XI0 vdd vss in<2> in<0> in<1> out<0> out<1> out<2> out<3> / 2x4decoder
XI2 in<2> inn<2> vdd vss / inv1
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    4x16decoder
* View Name:    schematic
************************************************************************

.SUBCKT 4x16decoder VDD VSS en in<0> in<1> in<2> in<3> out<0> out<1> out<2> 
+ out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11> out<12> 
+ out<13> out<14> out<15>
*.PININFO en:I in<0>:I in<1>:I in<2>:I in<3>:I out<0>:O out<1>:O out<2>:O 
*.PININFO out<3>:O out<4>:O out<5>:O out<6>:O out<7>:O out<8>:O out<9>:O 
*.PININFO out<10>:O out<11>:O out<12>:O out<13>:O out<14>:O out<15>:O VDD:B 
*.PININFO VSS:B
XI15 VDD VSS en in<2> in<3> b<0> b<1> b<2> b<3> / 2x4decoder
XI0 VDD VSS en in<0> in<1> c<0> c<1> c<2> c<3> / 2x4decoder
XI73 net173 out<15> VDD VSS / inv4
XI70 net174 out<14> VDD VSS / inv4
XI69 net175 out<13> VDD VSS / inv4
XI67 net176 out<12> VDD VSS / inv4
XI81 net092 out<11> VDD VSS / inv4
XI78 net097 out<10> VDD VSS / inv4
XI77 net179 out<9> VDD VSS / inv4
XI75 net180 out<8> VDD VSS / inv4
XI65 net0112 out<7> VDD VSS / inv4
XI62 net182 out<6> VDD VSS / inv4
XI61 net183 out<5> VDD VSS / inv4
XI59 net0127 out<4> VDD VSS / inv4
XI57 net185 out<3> VDD VSS / inv4
XI54 net0137 out<2> VDD VSS / inv4
XI53 net187 out<1> VDD VSS / inv4
XI51 net188 out<0> VDD VSS / inv4
XI8 c<2> b<2> net097 VDD VSS / nand
XI7 c<3> b<2> net092 VDD VSS / nand
XI6 c<3> b<1> net0112 VDD VSS / nand
XI5 c<2> b<1> net182 VDD VSS / nand
XI4 c<0> b<1> net0127 VDD VSS / nand
XI3 c<1> b<1> net183 VDD VSS / nand
XI2 c<3> b<0> net185 VDD VSS / nand
XI1 c<2> b<0> net0137 VDD VSS / nand
XI9 c<0> b<2> net180 VDD VSS / nand
XI10 c<1> b<2> net179 VDD VSS / nand
XI11 c<1> b<3> net175 VDD VSS / nand
XI12 c<0> b<3> net176 VDD VSS / nand
XI13 c<2> b<3> net174 VDD VSS / nand
XI14 c<3> b<3> net173 VDD VSS / nand
XI50 c<0> b<0> net188 VDD VSS / nand
XI52 c<1> b<0> net187 VDD VSS / nand
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    access_decoder
* View Name:    schematic
************************************************************************

.SUBCKT access_decoder a_col<0> a_col<1> a_row<0> a_row<1> a_row<2> a_row<3> 
+ a_row<4> a_row<5> a_row<6> col<0> col<1> col<2> col<3> en_acc_col en_acc_row 
+ group<0> group<1> group<2> group<3> group<4> group<5> group<6> group<7> 
+ row16<0> row16<1> row16<2> row16<3> row16<4> row16<5> row16<6> row16<7> 
+ row16<8> row16<9> row16<10> row16<11> row16<12> row16<13> row16<14> 
+ row16<15> vdd vss wrt wrtbuf
*.PININFO a_col<0>:I a_col<1>:I a_row<0>:I a_row<1>:I a_row<2>:I a_row<3>:I 
*.PININFO a_row<4>:I a_row<5>:I a_row<6>:I en_acc_col:I en_acc_row:I col<0>:O 
*.PININFO col<1>:O col<2>:O col<3>:O group<0>:O group<1>:O group<2>:O 
*.PININFO group<3>:O group<4>:O group<5>:O group<6>:O group<7>:O row16<0>:O 
*.PININFO row16<1>:O row16<2>:O row16<3>:O row16<4>:O row16<5>:O row16<6>:O 
*.PININFO row16<7>:O row16<8>:O row16<9>:O row16<10>:O row16<11>:O row16<12>:O 
*.PININFO row16<13>:O row16<14>:O row16<15>:O vdd:B vss:B wrt:B wrtbuf:B
XI0 a_row<0> a_row<1> a_row<2> group<0> group<1> group<2> group<3> group<4> 
+ group<5> group<6> group<7> vdd vss / 3x8decoder
XI1 vdd vss en_acc_row a_row<3> a_row<4> a_row<5> a_row<6> row16<0> row16<1> 
+ row16<2> row16<3> row16<4> row16<5> row16<6> row16<7> row16<8> row16<9> 
+ row16<10> row16<11> row16<12> row16<13> row16<14> row16<15> / 4x16decoder
XI2 vdd vss en_acc_col a_col<0> a_col<1> col<0> col<1> col<2> col<3> / 
+ 2x4decoder
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    master
* View Name:    schematic
************************************************************************

.SUBCKT master a<0> a<1> a<2> a<3> a<4> a<5> a<6> a<7> a<8> a_col<0> a_col<1> 
+ a_inbuf<0> a_inbuf<1> a_inbuf<2> a_inbuf<3> a_inbuf<4> a_read<0> a_read<1> 
+ a_read<2> a_read<3> a_row<0> a_row<1> a_row<2> a_row<3> a_row<4> a_row<5> 
+ a_row<6> clk clk_read clk_write comp en_acc_col en_acc_row eninbuf enread 
+ entime inbit model model_ read set set_ set_comp time<0> time<1> time<2> 
+ time<3> vdd vss wait wrt wrt_ wrtbuf wrtbuf_
*.PININFO a<0>:I a<1>:I a<2>:I a<3>:I a<4>:I a<5>:I a<6>:I a<7>:I a<8>:I clk:I 
*.PININFO comp:I inbit:I model:I read:I set:I wait:I wrt:I wrtbuf:I a_col<0>:O 
*.PININFO a_col<1>:O a_inbuf<0>:O a_inbuf<1>:O a_inbuf<2>:O a_inbuf<3>:O 
*.PININFO a_inbuf<4>:O a_read<0>:O a_read<1>:O a_read<2>:O a_read<3>:O 
*.PININFO a_row<0>:O a_row<1>:O a_row<2>:O a_row<3>:O a_row<4>:O a_row<5>:O 
*.PININFO a_row<6>:O clk_read:O clk_write:O en_acc_col:O en_acc_row:O 
*.PININFO eninbuf:O enread:O entime:O model_:O set_:O set_comp:O time<0>:O 
*.PININFO time<1>:O time<2>:O time<3>:O wrt_:O wrtbuf_:O vdd:B vss:B
XI102 net015 waitb vdd vss / inv2
XI114 net018 net049 vdd vss / inv2
XI113 net019 net018 vdd vss / inv2
XI116 net0100 net039 vdd vss / inv2
XI115 net016 net0100 vdd vss / inv2
XI46 net077 net074 vdd vss / inv2
XI7 net051 compb vdd vss / inv2
XI5 net050 setb vdd vss / inv2
XI13 net040 readb vdd vss / inv2
XI15 net039 inbitb vdd vss / inv2
XI2 net049 modelb vdd vss / inv2
XI17 net038 wrtbufb vdd vss / inv2
XI1<0> net054<0> ab<0> vdd vss / inv2
XI1<1> net054<1> ab<1> vdd vss / inv2
XI1<2> net054<2> ab<2> vdd vss / inv2
XI1<3> net054<3> ab<3> vdd vss / inv2
XI1<4> net054<4> ab<4> vdd vss / inv2
XI1<5> net054<5> ab<5> vdd vss / inv2
XI1<6> net054<6> ab<6> vdd vss / inv2
XI1<7> net054<7> ab<7> vdd vss / inv2
XI1<8> net054<8> ab<8> vdd vss / inv2
XI11 net053 wrtb vdd vss / inv2
XI101 wait net015 vdd vss / inv8
XI65<0> net084<0> a_row<0> vdd vss / inv8
XI65<1> net084<1> a_row<1> vdd vss / inv8
XI65<2> net084<2> a_row<2> vdd vss / inv8
XI65<3> net084<3> a_row<3> vdd vss / inv8
XI65<4> net084<4> a_row<4> vdd vss / inv8
XI65<5> net084<5> a_row<5> vdd vss / inv8
XI65<6> net084<6> a_row<6> vdd vss / inv8
XI70<0> net085<0> a_col<0> vdd vss / inv8
XI70<1> net085<1> a_col<1> vdd vss / inv8
XI72<0> net059<0> a_read<0> vdd vss / inv8
XI72<1> net059<1> a_read<1> vdd vss / inv8
XI72<2> net059<2> a_read<2> vdd vss / inv8
XI72<3> net059<3> a_read<3> vdd vss / inv8
XI68<0> net060<0> a_inbuf<0> vdd vss / inv8
XI68<1> net060<1> a_inbuf<1> vdd vss / inv8
XI68<2> net060<2> a_inbuf<2> vdd vss / inv8
XI68<3> net060<3> a_inbuf<3> vdd vss / inv8
XI68<4> net060<4> a_inbuf<4> vdd vss / inv8
XI59 net064 eninbuf vdd vss / inv8
XI58 net067 en_acc_col vdd vss / inv8
XI56 net068 en_acc_row vdd vss / inv8
XI53 net069 enread vdd vss / inv8
XI49 net070 set_comp vdd vss / inv8
XI43 net076 clk_write vdd vss / inv8
XI39 net062 clk_read vdd vss / inv8
XI31 net080 set_ vdd vss / inv8
XI30 net081 model_ vdd vss / inv8
XI0<0> a<0> net054<0> vdd vss / inv8
XI0<1> a<1> net054<1> vdd vss / inv8
XI0<2> a<2> net054<2> vdd vss / inv8
XI0<3> a<3> net054<3> vdd vss / inv8
XI0<4> a<4> net054<4> vdd vss / inv8
XI0<5> a<5> net054<5> vdd vss / inv8
XI0<6> a<6> net054<6> vdd vss / inv8
XI0<7> a<7> net054<7> vdd vss / inv8
XI0<8> a<8> net054<8> vdd vss / inv8
XI8 clk net052 vdd vss / inv8
XI9 net052 clkb vdd vss / inv8
XI6 comp net051 vdd vss / inv8
XI4 set net050 vdd vss / inv8
XI14 inbit net016 vdd vss / inv8
XI12 read net040 vdd vss / inv8
XI16 wrtbuf net038 vdd vss / inv8
XI26 net061 wrtbuf_ vdd vss / inv8
XI19 net06 wrt_ vdd vss / inv8
XI3 model net019 vdd vss / inv8
XI10 wrt net053 vdd vss / inv8
XI112 clkcharge net026 net022 vdd vss / nand
XI110 clkcharge net025 net023 vdd vss / nand
XI108 clkcharge net027 net024 vdd vss / nand
XI106 clkcharge net029 net028 vdd vss / nand
XI104 clkb net012 net097 vdd vss / nand
XI99 net0126 inbitb net0132 vdd vss / nand
XI96 compb modelb net0128 vdd vss / nand
XI93 net066 inbitn net065 vdd vss / nand
XI90 compb modelb net0122 vdd vss / nand
XI87 net0137 inbitb net0124 vdd vss / nand
XI84 compb modeln net0121 vdd vss / nand
XI81 net0131 inbitn net0120 vdd vss / nand
XI78 compb modeln net0136 vdd vss / nand
XI47 net074 clkb net075 vdd vss / nand
XI37 clkb readb net079 vdd vss / nand
XI20 clkb wrtbufb net014 vdd vss / nand
XI18 clkb wrtb net013 vdd vss / nand
XI111 net022 time<0> vdd vss / inv4
XI109 net023 time<1> vdd vss / inv4
XI107 net024 time<2> vdd vss / inv4
XI105 net028 time<3> vdd vss / inv4
XI103 net097 clkcharge vdd vss / inv4
XI98 net0132 net029 vdd vss / inv4
XI97 net0128 net0126 vdd vss / inv4
XI92 net065 net027 vdd vss / inv4
XI91 net0122 net066 vdd vss / inv4
XI86 net0124 net025 vdd vss / inv4
XI85 net0121 net0137 vdd vss / inv4
XI69<0> ab<7> net085<0> vdd vss / inv4
XI69<1> ab<8> net085<1> vdd vss / inv4
XI75 inbitb inbitn vdd vss / inv4
XI67<0> ab<0> net060<0> vdd vss / inv4
XI67<1> ab<1> net060<1> vdd vss / inv4
XI67<2> ab<2> net060<2> vdd vss / inv4
XI67<3> ab<3> net060<3> vdd vss / inv4
XI67<4> ab<4> net060<4> vdd vss / inv4
XI71<0> ab<0> net059<0> vdd vss / inv4
XI71<1> ab<1> net059<1> vdd vss / inv4
XI71<2> ab<2> net059<2> vdd vss / inv4
XI71<3> ab<3> net059<3> vdd vss / inv4
XI80 net0120 net026 vdd vss / inv4
XI79 net0136 net0131 vdd vss / inv4
XI66<0> ab<0> net084<0> vdd vss / inv4
XI66<1> ab<1> net084<1> vdd vss / inv4
XI66<2> ab<2> net084<2> vdd vss / inv4
XI66<3> ab<3> net084<3> vdd vss / inv4
XI66<4> ab<4> net084<4> vdd vss / inv4
XI66<5> ab<5> net084<5> vdd vss / inv4
XI66<6> ab<6> net084<6> vdd vss / inv4
XI119 net095 net012 vdd vss / inv4
XI60 net061 net064 vdd vss / inv4
XI57 net06 net067 vdd vss / inv4
XI55 net06 net068 vdd vss / inv4
XI54 net062 net069 vdd vss / inv4
XI52 net072 net071 vdd vss / inv4
XI50 net071 net070 vdd vss / inv4
XI48 net075 net073 vdd vss / inv4
XI44 net073 net076 vdd vss / inv4
XI38 net079 net078 vdd vss / inv4
XI40 net078 net062 vdd vss / inv4
XI117 net071 entime vdd vss / inv4
XI82 modelb modeln vdd vss / inv4
XI32 setb net080 vdd vss / inv4
XI29 modelb net081 vdd vss / inv4
XI25 net011 net06 vdd vss / inv4
XI28 net082 net061 vdd vss / inv4
XI27 net014 net082 vdd vss / inv4
XI22 net013 net011 vdd vss / inv4
XI118 waitb setb net095 vdd vss / nor
XI51 setb compb net072 vdd vss / nor
XI45 wrtb wrtbufb net077 vdd vss / nor
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    inputsinglecell
* View Name:    schematic
************************************************************************

.SUBCKT inputsinglecell bl<0> bl<1> bl<2> bl<3> q<0> q<1> q<2> q<3> sl<0> 
+ sl<1> sl<2> sl<3> vdd vss wl
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I sl<0>:I sl<1>:I sl<2>:I sl<3>:I wl:I 
*.PININFO q<0>:O q<1>:O q<2>:O q<3>:O vdd:B vss:B
XI3 bl<3> q<3> net18 sl<3> vdd vss wl / cell_SRAM
XI2 bl<0> q<0> net19 sl<0> vdd vss wl / cell_SRAM
XI1 bl<2> q<2> net20 sl<2> vdd vss wl / cell_SRAM
XI0 bl<1> q<1> net21 sl<1> vdd vss wl / cell_SRAM
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    inputcell
* View Name:    schematic
************************************************************************

.SUBCKT inputcell bl<0> bl<1> bl<2> bl<3> q0<0> q0<1> q0<2> q0<3> q0<4> q0<5> 
+ q0<6> q0<7> q0<8> q0<9> q0<10> q0<11> q0<12> q0<13> q0<14> q0<15> q0<16> 
+ q0<17> q0<18> q0<19> q0<20> q0<21> q0<22> q0<23> q0<24> q0<25> q0<26> q0<27> 
+ q0<28> q0<29> q0<30> q0<31> q1<0> q1<1> q1<2> q1<3> q1<4> q1<5> q1<6> q1<7> 
+ q1<8> q1<9> q1<10> q1<11> q1<12> q1<13> q1<14> q1<15> q1<16> q1<17> q1<18> 
+ q1<19> q1<20> q1<21> q1<22> q1<23> q1<24> q1<25> q1<26> q1<27> q1<28> q1<29> 
+ q1<30> q1<31> q2<0> q2<1> q2<2> q2<3> q2<4> q2<5> q2<6> q2<7> q2<8> q2<9> 
+ q2<10> q2<11> q2<12> q2<13> q2<14> q2<15> q2<16> q2<17> q2<18> q2<19> q2<20> 
+ q2<21> q2<22> q2<23> q2<24> q2<25> q2<26> q2<27> q2<28> q2<29> q2<30> q2<31> 
+ q3<0> q3<1> q3<2> q3<3> q3<4> q3<5> q3<6> q3<7> q3<8> q3<9> q3<10> q3<11> 
+ q3<12> q3<13> q3<14> q3<15> q3<16> q3<17> q3<18> q3<19> q3<20> q3<21> q3<22> 
+ q3<23> q3<24> q3<25> q3<26> q3<27> q3<28> q3<29> q3<30> q3<31> sl<0> sl<1> 
+ sl<2> sl<3> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> 
+ wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> 
+ wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> 
+ wl<31>
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I sl<0>:I sl<1>:I sl<2>:I sl<3>:I 
*.PININFO vdd:I vss:I wl<0>:I wl<1>:I wl<2>:I wl<3>:I wl<4>:I wl<5>:I wl<6>:I 
*.PININFO wl<7>:I wl<8>:I wl<9>:I wl<10>:I wl<11>:I wl<12>:I wl<13>:I wl<14>:I 
*.PININFO wl<15>:I wl<16>:I wl<17>:I wl<18>:I wl<19>:I wl<20>:I wl<21>:I 
*.PININFO wl<22>:I wl<23>:I wl<24>:I wl<25>:I wl<26>:I wl<27>:I wl<28>:I 
*.PININFO wl<29>:I wl<30>:I wl<31>:I q0<0>:O q0<1>:O q0<2>:O q0<3>:O q0<4>:O 
*.PININFO q0<5>:O q0<6>:O q0<7>:O q0<8>:O q0<9>:O q0<10>:O q0<11>:O q0<12>:O 
*.PININFO q0<13>:O q0<14>:O q0<15>:O q0<16>:O q0<17>:O q0<18>:O q0<19>:O 
*.PININFO q0<20>:O q0<21>:O q0<22>:O q0<23>:O q0<24>:O q0<25>:O q0<26>:O 
*.PININFO q0<27>:O q0<28>:O q0<29>:O q0<30>:O q0<31>:O q1<0>:O q1<1>:O q1<2>:O 
*.PININFO q1<3>:O q1<4>:O q1<5>:O q1<6>:O q1<7>:O q1<8>:O q1<9>:O q1<10>:O 
*.PININFO q1<11>:O q1<12>:O q1<13>:O q1<14>:O q1<15>:O q1<16>:O q1<17>:O 
*.PININFO q1<18>:O q1<19>:O q1<20>:O q1<21>:O q1<22>:O q1<23>:O q1<24>:O 
*.PININFO q1<25>:O q1<26>:O q1<27>:O q1<28>:O q1<29>:O q1<30>:O q1<31>:O 
*.PININFO q2<0>:O q2<1>:O q2<2>:O q2<3>:O q2<4>:O q2<5>:O q2<6>:O q2<7>:O 
*.PININFO q2<8>:O q2<9>:O q2<10>:O q2<11>:O q2<12>:O q2<13>:O q2<14>:O 
*.PININFO q2<15>:O q2<16>:O q2<17>:O q2<18>:O q2<19>:O q2<20>:O q2<21>:O 
*.PININFO q2<22>:O q2<23>:O q2<24>:O q2<25>:O q2<26>:O q2<27>:O q2<28>:O 
*.PININFO q2<29>:O q2<30>:O q2<31>:O q3<0>:O q3<1>:O q3<2>:O q3<3>:O q3<4>:O 
*.PININFO q3<5>:O q3<6>:O q3<7>:O q3<8>:O q3<9>:O q3<10>:O q3<11>:O q3<12>:O 
*.PININFO q3<13>:O q3<14>:O q3<15>:O q3<16>:O q3<17>:O q3<18>:O q3<19>:O 
*.PININFO q3<20>:O q3<21>:O q3<22>:O q3<23>:O q3<24>:O q3<25>:O q3<26>:O 
*.PININFO q3<27>:O q3<28>:O q3<29>:O q3<30>:O q3<31>:O
XI167 bl<0> bl<1> bl<2> bl<3> q0<0> q1<0> q2<0> q3<0> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<0> / inputsinglecell
XI168 bl<0> bl<1> bl<2> bl<3> q0<1> q1<1> q2<1> q3<1> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<1> / inputsinglecell
XI169 bl<0> bl<1> bl<2> bl<3> q0<2> q1<2> q2<2> q3<2> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<2> / inputsinglecell
XI170 bl<0> bl<1> bl<2> bl<3> q0<3> q1<3> q2<3> q3<3> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<3> / inputsinglecell
XI171 bl<0> bl<1> bl<2> bl<3> q0<4> q1<4> q2<4> q3<4> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<4> / inputsinglecell
XI172 bl<0> bl<1> bl<2> bl<3> q0<5> q1<5> q2<5> q3<5> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<5> / inputsinglecell
XI173 bl<0> bl<1> bl<2> bl<3> q0<6> q1<6> q2<6> q3<6> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<6> / inputsinglecell
XI174 bl<0> bl<1> bl<2> bl<3> q0<7> q1<7> q2<7> q3<7> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<7> / inputsinglecell
XI175 bl<0> bl<1> bl<2> bl<3> q0<8> q1<8> q2<8> q3<8> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<8> / inputsinglecell
XI176 bl<0> bl<1> bl<2> bl<3> q0<9> q1<9> q2<9> q3<9> sl<0> sl<1> sl<2> sl<3> 
+ vdd vss wl<9> / inputsinglecell
XI177 bl<0> bl<1> bl<2> bl<3> q0<10> q1<10> q2<10> q3<10> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<10> / inputsinglecell
XI178 bl<0> bl<1> bl<2> bl<3> q0<11> q1<11> q2<11> q3<11> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<11> / inputsinglecell
XI179 bl<0> bl<1> bl<2> bl<3> q0<12> q1<12> q2<12> q3<12> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<12> / inputsinglecell
XI180 bl<0> bl<1> bl<2> bl<3> q0<13> q1<13> q2<13> q3<13> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<13> / inputsinglecell
XI181 bl<0> bl<1> bl<2> bl<3> q0<14> q1<14> q2<14> q3<14> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<14> / inputsinglecell
XI182 bl<0> bl<1> bl<2> bl<3> q0<15> q1<15> q2<15> q3<15> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<15> / inputsinglecell
XI183 bl<0> bl<1> bl<2> bl<3> q0<16> q1<16> q2<16> q3<16> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<16> / inputsinglecell
XI184 bl<0> bl<1> bl<2> bl<3> q0<17> q1<17> q2<17> q3<17> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<17> / inputsinglecell
XI185 bl<0> bl<1> bl<2> bl<3> q0<18> q1<18> q2<18> q3<18> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<18> / inputsinglecell
XI186 bl<0> bl<1> bl<2> bl<3> q0<19> q1<19> q2<19> q3<19> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<19> / inputsinglecell
XI187 bl<0> bl<1> bl<2> bl<3> q0<20> q1<20> q2<20> q3<20> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<20> / inputsinglecell
XI188 bl<0> bl<1> bl<2> bl<3> q0<21> q1<21> q2<21> q3<21> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<21> / inputsinglecell
XI189 bl<0> bl<1> bl<2> bl<3> q0<22> q1<22> q2<22> q3<22> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<22> / inputsinglecell
XI190 bl<0> bl<1> bl<2> bl<3> q0<23> q1<23> q2<23> q3<23> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<23> / inputsinglecell
XI191 bl<0> bl<1> bl<2> bl<3> q0<24> q1<24> q2<24> q3<24> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<24> / inputsinglecell
XI192 bl<0> bl<1> bl<2> bl<3> q0<25> q1<25> q2<25> q3<25> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<25> / inputsinglecell
XI193 bl<0> bl<1> bl<2> bl<3> q0<26> q1<26> q2<26> q3<26> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<26> / inputsinglecell
XI194 bl<0> bl<1> bl<2> bl<3> q0<27> q1<27> q2<27> q3<27> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<27> / inputsinglecell
XI195 bl<0> bl<1> bl<2> bl<3> q0<28> q1<28> q2<28> q3<28> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<28> / inputsinglecell
XI196 bl<0> bl<1> bl<2> bl<3> q0<29> q1<29> q2<29> q3<29> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<29> / inputsinglecell
XI197 bl<0> bl<1> bl<2> bl<3> q0<30> q1<30> q2<30> q3<30> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<30> / inputsinglecell
XI198 bl<0> bl<1> bl<2> bl<3> q0<31> q1<31> q2<31> q3<31> sl<0> sl<1> sl<2> 
+ sl<3> vdd vss wl<31> / inputsinglecell
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    inputbuffer
* View Name:    schematic
************************************************************************

.SUBCKT inputbuffer bl<0> bl<1> bl<2> bl<3> bl<4> bl<5> bl<6> bl<7> bl<8> 
+ bl<9> bl<10> bl<11> bl<12> bl<13> bl<14> bl<15> q0<0> q0<1> q0<2> q0<3> 
+ q0<4> q0<5> q0<6> q0<7> q0<8> q0<9> q0<10> q0<11> q0<12> q0<13> q0<14> 
+ q0<15> q0<16> q0<17> q0<18> q0<19> q0<20> q0<21> q0<22> q0<23> q0<24> q0<25> 
+ q0<26> q0<27> q0<28> q0<29> q0<30> q0<31> q0<32> q0<33> q0<34> q0<35> q0<36> 
+ q0<37> q0<38> q0<39> q0<40> q0<41> q0<42> q0<43> q0<44> q0<45> q0<46> q0<47> 
+ q0<48> q0<49> q0<50> q0<51> q0<52> q0<53> q0<54> q0<55> q0<56> q0<57> q0<58> 
+ q0<59> q0<60> q0<61> q0<62> q0<63> q0<64> q0<65> q0<66> q0<67> q0<68> q0<69> 
+ q0<70> q0<71> q0<72> q0<73> q0<74> q0<75> q0<76> q0<77> q0<78> q0<79> q0<80> 
+ q0<81> q0<82> q0<83> q0<84> q0<85> q0<86> q0<87> q0<88> q0<89> q0<90> q0<91> 
+ q0<92> q0<93> q0<94> q0<95> q0<96> q0<97> q0<98> q0<99> q0<100> q0<101> 
+ q0<102> q0<103> q0<104> q0<105> q0<106> q0<107> q0<108> q0<109> q0<110> 
+ q0<111> q0<112> q0<113> q0<114> q0<115> q0<116> q0<117> q0<118> q0<119> 
+ q0<120> q0<121> q0<122> q0<123> q0<124> q0<125> q0<126> q0<127> q1<0> q1<1> 
+ q1<2> q1<3> q1<4> q1<5> q1<6> q1<7> q1<8> q1<9> q1<10> q1<11> q1<12> q1<13> 
+ q1<14> q1<15> q1<16> q1<17> q1<18> q1<19> q1<20> q1<21> q1<22> q1<23> q1<24> 
+ q1<25> q1<26> q1<27> q1<28> q1<29> q1<30> q1<31> q1<32> q1<33> q1<34> q1<35> 
+ q1<36> q1<37> q1<38> q1<39> q1<40> q1<41> q1<42> q1<43> q1<44> q1<45> q1<46> 
+ q1<47> q1<48> q1<49> q1<50> q1<51> q1<52> q1<53> q1<54> q1<55> q1<56> q1<57> 
+ q1<58> q1<59> q1<60> q1<61> q1<62> q1<63> q1<64> q1<65> q1<66> q1<67> q1<68> 
+ q1<69> q1<70> q1<71> q1<72> q1<73> q1<74> q1<75> q1<76> q1<77> q1<78> q1<79> 
+ q1<80> q1<81> q1<82> q1<83> q1<84> q1<85> q1<86> q1<87> q1<88> q1<89> q1<90> 
+ q1<91> q1<92> q1<93> q1<94> q1<95> q1<96> q1<97> q1<98> q1<99> q1<100> 
+ q1<101> q1<102> q1<103> q1<104> q1<105> q1<106> q1<107> q1<108> q1<109> 
+ q1<110> q1<111> q1<112> q1<113> q1<114> q1<115> q1<116> q1<117> q1<118> 
+ q1<119> q1<120> q1<121> q1<122> q1<123> q1<124> q1<125> q1<126> q1<127> 
+ q2<0> q2<1> q2<2> q2<3> q2<4> q2<5> q2<6> q2<7> q2<8> q2<9> q2<10> q2<11> 
+ q2<12> q2<13> q2<14> q2<15> q2<16> q2<17> q2<18> q2<19> q2<20> q2<21> q2<22> 
+ q2<23> q2<24> q2<25> q2<26> q2<27> q2<28> q2<29> q2<30> q2<31> q2<32> q2<33> 
+ q2<34> q2<35> q2<36> q2<37> q2<38> q2<39> q2<40> q2<41> q2<42> q2<43> q2<44> 
+ q2<45> q2<46> q2<47> q2<48> q2<49> q2<50> q2<51> q2<52> q2<53> q2<54> q2<55> 
+ q2<56> q2<57> q2<58> q2<59> q2<60> q2<61> q2<62> q2<63> q2<64> q2<65> q2<66> 
+ q2<67> q2<68> q2<69> q2<70> q2<71> q2<72> q2<73> q2<74> q2<75> q2<76> q2<77> 
+ q2<78> q2<79> q2<80> q2<81> q2<82> q2<83> q2<84> q2<85> q2<86> q2<87> q2<88> 
+ q2<89> q2<90> q2<91> q2<92> q2<93> q2<94> q2<95> q2<96> q2<97> q2<98> q2<99> 
+ q2<100> q2<101> q2<102> q2<103> q2<104> q2<105> q2<106> q2<107> q2<108> 
+ q2<109> q2<110> q2<111> q2<112> q2<113> q2<114> q2<115> q2<116> q2<117> 
+ q2<118> q2<119> q2<120> q2<121> q2<122> q2<123> q2<124> q2<125> q2<126> 
+ q2<127> q3<0> q3<1> q3<2> q3<3> q3<4> q3<5> q3<6> q3<7> q3<8> q3<9> q3<10> 
+ q3<11> q3<12> q3<13> q3<14> q3<15> q3<16> q3<17> q3<18> q3<19> q3<20> q3<21> 
+ q3<22> q3<23> q3<24> q3<25> q3<26> q3<27> q3<28> q3<29> q3<30> q3<31> q3<32> 
+ q3<33> q3<34> q3<35> q3<36> q3<37> q3<38> q3<39> q3<40> q3<41> q3<42> q3<43> 
+ q3<44> q3<45> q3<46> q3<47> q3<48> q3<49> q3<50> q3<51> q3<52> q3<53> q3<54> 
+ q3<55> q3<56> q3<57> q3<58> q3<59> q3<60> q3<61> q3<62> q3<63> q3<64> q3<65> 
+ q3<66> q3<67> q3<68> q3<69> q3<70> q3<71> q3<72> q3<73> q3<74> q3<75> q3<76> 
+ q3<77> q3<78> q3<79> q3<80> q3<81> q3<82> q3<83> q3<84> q3<85> q3<86> q3<87> 
+ q3<88> q3<89> q3<90> q3<91> q3<92> q3<93> q3<94> q3<95> q3<96> q3<97> q3<98> 
+ q3<99> q3<100> q3<101> q3<102> q3<103> q3<104> q3<105> q3<106> q3<107> 
+ q3<108> q3<109> q3<110> q3<111> q3<112> q3<113> q3<114> q3<115> q3<116> 
+ q3<117> q3<118> q3<119> q3<120> q3<121> q3<122> q3<123> q3<124> q3<125> 
+ q3<126> q3<127> sl<0> sl<1> sl<2> sl<3> sl<4> sl<5> sl<6> sl<7> sl<8> sl<9> 
+ sl<10> sl<11> sl<12> sl<13> sl<14> sl<15> vdd vss wl<0> wl<1> wl<2> wl<3> 
+ wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> 
+ wl<15> wl<16> wl<17> wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> 
+ wl<26> wl<27> wl<28> wl<29> wl<30> wl<31>
*.PININFO bl<0>:I bl<1>:I bl<2>:I bl<3>:I bl<4>:I bl<5>:I bl<6>:I bl<7>:I 
*.PININFO bl<8>:I bl<9>:I bl<10>:I bl<11>:I bl<12>:I bl<13>:I bl<14>:I 
*.PININFO bl<15>:I sl<0>:I sl<1>:I sl<2>:I sl<3>:I sl<4>:I sl<5>:I sl<6>:I 
*.PININFO sl<7>:I sl<8>:I sl<9>:I sl<10>:I sl<11>:I sl<12>:I sl<13>:I sl<14>:I 
*.PININFO sl<15>:I wl<0>:I wl<1>:I wl<2>:I wl<3>:I wl<4>:I wl<5>:I wl<6>:I 
*.PININFO wl<7>:I wl<8>:I wl<9>:I wl<10>:I wl<11>:I wl<12>:I wl<13>:I wl<14>:I 
*.PININFO wl<15>:I wl<16>:I wl<17>:I wl<18>:I wl<19>:I wl<20>:I wl<21>:I 
*.PININFO wl<22>:I wl<23>:I wl<24>:I wl<25>:I wl<26>:I wl<27>:I wl<28>:I 
*.PININFO wl<29>:I wl<30>:I wl<31>:I q0<0>:O q0<1>:O q0<2>:O q0<3>:O q0<4>:O 
*.PININFO q0<5>:O q0<6>:O q0<7>:O q0<8>:O q0<9>:O q0<10>:O q0<11>:O q0<12>:O 
*.PININFO q0<13>:O q0<14>:O q0<15>:O q0<16>:O q0<17>:O q0<18>:O q0<19>:O 
*.PININFO q0<20>:O q0<21>:O q0<22>:O q0<23>:O q0<24>:O q0<25>:O q0<26>:O 
*.PININFO q0<27>:O q0<28>:O q0<29>:O q0<30>:O q0<31>:O q0<32>:O q0<33>:O 
*.PININFO q0<34>:O q0<35>:O q0<36>:O q0<37>:O q0<38>:O q0<39>:O q0<40>:O 
*.PININFO q0<41>:O q0<42>:O q0<43>:O q0<44>:O q0<45>:O q0<46>:O q0<47>:O 
*.PININFO q0<48>:O q0<49>:O q0<50>:O q0<51>:O q0<52>:O q0<53>:O q0<54>:O 
*.PININFO q0<55>:O q0<56>:O q0<57>:O q0<58>:O q0<59>:O q0<60>:O q0<61>:O 
*.PININFO q0<62>:O q0<63>:O q0<64>:O q0<65>:O q0<66>:O q0<67>:O q0<68>:O 
*.PININFO q0<69>:O q0<70>:O q0<71>:O q0<72>:O q0<73>:O q0<74>:O q0<75>:O 
*.PININFO q0<76>:O q0<77>:O q0<78>:O q0<79>:O q0<80>:O q0<81>:O q0<82>:O 
*.PININFO q0<83>:O q0<84>:O q0<85>:O q0<86>:O q0<87>:O q0<88>:O q0<89>:O 
*.PININFO q0<90>:O q0<91>:O q0<92>:O q0<93>:O q0<94>:O q0<95>:O q0<96>:O 
*.PININFO q0<97>:O q0<98>:O q0<99>:O q0<100>:O q0<101>:O q0<102>:O q0<103>:O 
*.PININFO q0<104>:O q0<105>:O q0<106>:O q0<107>:O q0<108>:O q0<109>:O 
*.PININFO q0<110>:O q0<111>:O q0<112>:O q0<113>:O q0<114>:O q0<115>:O 
*.PININFO q0<116>:O q0<117>:O q0<118>:O q0<119>:O q0<120>:O q0<121>:O 
*.PININFO q0<122>:O q0<123>:O q0<124>:O q0<125>:O q0<126>:O q0<127>:O q1<0>:O 
*.PININFO q1<1>:O q1<2>:O q1<3>:O q1<4>:O q1<5>:O q1<6>:O q1<7>:O q1<8>:O 
*.PININFO q1<9>:O q1<10>:O q1<11>:O q1<12>:O q1<13>:O q1<14>:O q1<15>:O 
*.PININFO q1<16>:O q1<17>:O q1<18>:O q1<19>:O q1<20>:O q1<21>:O q1<22>:O 
*.PININFO q1<23>:O q1<24>:O q1<25>:O q1<26>:O q1<27>:O q1<28>:O q1<29>:O 
*.PININFO q1<30>:O q1<31>:O q1<32>:O q1<33>:O q1<34>:O q1<35>:O q1<36>:O 
*.PININFO q1<37>:O q1<38>:O q1<39>:O q1<40>:O q1<41>:O q1<42>:O q1<43>:O 
*.PININFO q1<44>:O q1<45>:O q1<46>:O q1<47>:O q1<48>:O q1<49>:O q1<50>:O 
*.PININFO q1<51>:O q1<52>:O q1<53>:O q1<54>:O q1<55>:O q1<56>:O q1<57>:O 
*.PININFO q1<58>:O q1<59>:O q1<60>:O q1<61>:O q1<62>:O q1<63>:O q1<64>:O 
*.PININFO q1<65>:O q1<66>:O q1<67>:O q1<68>:O q1<69>:O q1<70>:O q1<71>:O 
*.PININFO q1<72>:O q1<73>:O q1<74>:O q1<75>:O q1<76>:O q1<77>:O q1<78>:O 
*.PININFO q1<79>:O q1<80>:O q1<81>:O q1<82>:O q1<83>:O q1<84>:O q1<85>:O 
*.PININFO q1<86>:O q1<87>:O q1<88>:O q1<89>:O q1<90>:O q1<91>:O q1<92>:O 
*.PININFO q1<93>:O q1<94>:O q1<95>:O q1<96>:O q1<97>:O q1<98>:O q1<99>:O 
*.PININFO q1<100>:O q1<101>:O q1<102>:O q1<103>:O q1<104>:O q1<105>:O 
*.PININFO q1<106>:O q1<107>:O q1<108>:O q1<109>:O q1<110>:O q1<111>:O 
*.PININFO q1<112>:O q1<113>:O q1<114>:O q1<115>:O q1<116>:O q1<117>:O 
*.PININFO q1<118>:O q1<119>:O q1<120>:O q1<121>:O q1<122>:O q1<123>:O 
*.PININFO q1<124>:O q1<125>:O q1<126>:O q1<127>:O q2<0>:O q2<1>:O q2<2>:O 
*.PININFO q2<3>:O q2<4>:O q2<5>:O q2<6>:O q2<7>:O q2<8>:O q2<9>:O q2<10>:O 
*.PININFO q2<11>:O q2<12>:O q2<13>:O q2<14>:O q2<15>:O q2<16>:O q2<17>:O 
*.PININFO q2<18>:O q2<19>:O q2<20>:O q2<21>:O q2<22>:O q2<23>:O q2<24>:O 
*.PININFO q2<25>:O q2<26>:O q2<27>:O q2<28>:O q2<29>:O q2<30>:O q2<31>:O 
*.PININFO q2<32>:O q2<33>:O q2<34>:O q2<35>:O q2<36>:O q2<37>:O q2<38>:O 
*.PININFO q2<39>:O q2<40>:O q2<41>:O q2<42>:O q2<43>:O q2<44>:O q2<45>:O 
*.PININFO q2<46>:O q2<47>:O q2<48>:O q2<49>:O q2<50>:O q2<51>:O q2<52>:O 
*.PININFO q2<53>:O q2<54>:O q2<55>:O q2<56>:O q2<57>:O q2<58>:O q2<59>:O 
*.PININFO q2<60>:O q2<61>:O q2<62>:O q2<63>:O q2<64>:O q2<65>:O q2<66>:O 
*.PININFO q2<67>:O q2<68>:O q2<69>:O q2<70>:O q2<71>:O q2<72>:O q2<73>:O 
*.PININFO q2<74>:O q2<75>:O q2<76>:O q2<77>:O q2<78>:O q2<79>:O q2<80>:O 
*.PININFO q2<81>:O q2<82>:O q2<83>:O q2<84>:O q2<85>:O q2<86>:O q2<87>:O 
*.PININFO q2<88>:O q2<89>:O q2<90>:O q2<91>:O q2<92>:O q2<93>:O q2<94>:O 
*.PININFO q2<95>:O q2<96>:O q2<97>:O q2<98>:O q2<99>:O q2<100>:O q2<101>:O 
*.PININFO q2<102>:O q2<103>:O q2<104>:O q2<105>:O q2<106>:O q2<107>:O 
*.PININFO q2<108>:O q2<109>:O q2<110>:O q2<111>:O q2<112>:O q2<113>:O 
*.PININFO q2<114>:O q2<115>:O q2<116>:O q2<117>:O q2<118>:O q2<119>:O 
*.PININFO q2<120>:O q2<121>:O q2<122>:O q2<123>:O q2<124>:O q2<125>:O 
*.PININFO q2<126>:O q2<127>:O q3<0>:O q3<1>:O q3<2>:O q3<3>:O q3<4>:O q3<5>:O 
*.PININFO q3<6>:O q3<7>:O q3<8>:O q3<9>:O q3<10>:O q3<11>:O q3<12>:O q3<13>:O 
*.PININFO q3<14>:O q3<15>:O q3<16>:O q3<17>:O q3<18>:O q3<19>:O q3<20>:O 
*.PININFO q3<21>:O q3<22>:O q3<23>:O q3<24>:O q3<25>:O q3<26>:O q3<27>:O 
*.PININFO q3<28>:O q3<29>:O q3<30>:O q3<31>:O q3<32>:O q3<33>:O q3<34>:O 
*.PININFO q3<35>:O q3<36>:O q3<37>:O q3<38>:O q3<39>:O q3<40>:O q3<41>:O 
*.PININFO q3<42>:O q3<43>:O q3<44>:O q3<45>:O q3<46>:O q3<47>:O q3<48>:O 
*.PININFO q3<49>:O q3<50>:O q3<51>:O q3<52>:O q3<53>:O q3<54>:O q3<55>:O 
*.PININFO q3<56>:O q3<57>:O q3<58>:O q3<59>:O q3<60>:O q3<61>:O q3<62>:O 
*.PININFO q3<63>:O q3<64>:O q3<65>:O q3<66>:O q3<67>:O q3<68>:O q3<69>:O 
*.PININFO q3<70>:O q3<71>:O q3<72>:O q3<73>:O q3<74>:O q3<75>:O q3<76>:O 
*.PININFO q3<77>:O q3<78>:O q3<79>:O q3<80>:O q3<81>:O q3<82>:O q3<83>:O 
*.PININFO q3<84>:O q3<85>:O q3<86>:O q3<87>:O q3<88>:O q3<89>:O q3<90>:O 
*.PININFO q3<91>:O q3<92>:O q3<93>:O q3<94>:O q3<95>:O q3<96>:O q3<97>:O 
*.PININFO q3<98>:O q3<99>:O q3<100>:O q3<101>:O q3<102>:O q3<103>:O q3<104>:O 
*.PININFO q3<105>:O q3<106>:O q3<107>:O q3<108>:O q3<109>:O q3<110>:O 
*.PININFO q3<111>:O q3<112>:O q3<113>:O q3<114>:O q3<115>:O q3<116>:O 
*.PININFO q3<117>:O q3<118>:O q3<119>:O q3<120>:O q3<121>:O q3<122>:O 
*.PININFO q3<123>:O q3<124>:O q3<125>:O q3<126>:O q3<127>:O vdd:B vss:B
XI4 bl<12> bl<13> bl<14> bl<15> q0<96> q0<97> q0<98> q0<99> q0<100> q0<101> 
+ q0<102> q0<103> q0<104> q0<105> q0<106> q0<107> q0<108> q0<109> q0<110> 
+ q0<111> q0<112> q0<113> q0<114> q0<115> q0<116> q0<117> q0<118> q0<119> 
+ q0<120> q0<121> q0<122> q0<123> q0<124> q0<125> q0<126> q0<127> q1<96> 
+ q1<97> q1<98> q1<99> q1<100> q1<101> q1<102> q1<103> q1<104> q1<105> q1<106> 
+ q1<107> q1<108> q1<109> q1<110> q1<111> q1<112> q1<113> q1<114> q1<115> 
+ q1<116> q1<117> q1<118> q1<119> q1<120> q1<121> q1<122> q1<123> q1<124> 
+ q1<125> q1<126> q1<127> q2<96> q2<97> q2<98> q2<99> q2<100> q2<101> q2<102> 
+ q2<103> q2<104> q2<105> q2<106> q2<107> q2<108> q2<109> q2<110> q2<111> 
+ q2<112> q2<113> q2<114> q2<115> q2<116> q2<117> q2<118> q2<119> q2<120> 
+ q2<121> q2<122> q2<123> q2<124> q2<125> q2<126> q2<127> q3<96> q3<97> q3<98> 
+ q3<99> q3<100> q3<101> q3<102> q3<103> q3<104> q3<105> q3<106> q3<107> 
+ q3<108> q3<109> q3<110> q3<111> q3<112> q3<113> q3<114> q3<115> q3<116> 
+ q3<117> q3<118> q3<119> q3<120> q3<121> q3<122> q3<123> q3<124> q3<125> 
+ q3<126> q3<127> sl<12> sl<13> sl<14> sl<15> vdd vss wl<0> wl<1> wl<2> wl<3> 
+ wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> 
+ wl<15> wl<16> wl<17> wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> 
+ wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> / inputcell
XI3 bl<8> bl<9> bl<10> bl<11> q0<64> q0<65> q0<66> q0<67> q0<68> q0<69> q0<70> 
+ q0<71> q0<72> q0<73> q0<74> q0<75> q0<76> q0<77> q0<78> q0<79> q0<80> q0<81> 
+ q0<82> q0<83> q0<84> q0<85> q0<86> q0<87> q0<88> q0<89> q0<90> q0<91> q0<92> 
+ q0<93> q0<94> q0<95> q1<64> q1<65> q1<66> q1<67> q1<68> q1<69> q1<70> q1<71> 
+ q1<72> q1<73> q1<74> q1<75> q1<76> q1<77> q1<78> q1<79> q1<80> q1<81> q1<82> 
+ q1<83> q1<84> q1<85> q1<86> q1<87> q1<88> q1<89> q1<90> q1<91> q1<92> q1<93> 
+ q1<94> q1<95> q2<64> q2<65> q2<66> q2<67> q2<68> q2<69> q2<70> q2<71> q2<72> 
+ q2<73> q2<74> q2<75> q2<76> q2<77> q2<78> q2<79> q2<80> q2<81> q2<82> q2<83> 
+ q2<84> q2<85> q2<86> q2<87> q2<88> q2<89> q2<90> q2<91> q2<92> q2<93> q2<94> 
+ q2<95> q3<64> q3<65> q3<66> q3<67> q3<68> q3<69> q3<70> q3<71> q3<72> q3<73> 
+ q3<74> q3<75> q3<76> q3<77> q3<78> q3<79> q3<80> q3<81> q3<82> q3<83> q3<84> 
+ q3<85> q3<86> q3<87> q3<88> q3<89> q3<90> q3<91> q3<92> q3<93> q3<94> q3<95> 
+ sl<8> sl<9> sl<10> sl<11> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> 
+ wl<7> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> 
+ wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> 
+ wl<29> wl<30> wl<31> / inputcell
XI2 bl<4> bl<5> bl<6> bl<7> q0<32> q0<33> q0<34> q0<35> q0<36> q0<37> q0<38> 
+ q0<39> q0<40> q0<41> q0<42> q0<43> q0<44> q0<45> q0<46> q0<47> q0<48> q0<49> 
+ q0<50> q0<51> q0<52> q0<53> q0<54> q0<55> q0<56> q0<57> q0<58> q0<59> q0<60> 
+ q0<61> q0<62> q0<63> q1<32> q1<33> q1<34> q1<35> q1<36> q1<37> q1<38> q1<39> 
+ q1<40> q1<41> q1<42> q1<43> q1<44> q1<45> q1<46> q1<47> q1<48> q1<49> q1<50> 
+ q1<51> q1<52> q1<53> q1<54> q1<55> q1<56> q1<57> q1<58> q1<59> q1<60> q1<61> 
+ q1<62> q1<63> q2<32> q2<33> q2<34> q2<35> q2<36> q2<37> q2<38> q2<39> q2<40> 
+ q2<41> q2<42> q2<43> q2<44> q2<45> q2<46> q2<47> q2<48> q2<49> q2<50> q2<51> 
+ q2<52> q2<53> q2<54> q2<55> q2<56> q2<57> q2<58> q2<59> q2<60> q2<61> q2<62> 
+ q2<63> q3<32> q3<33> q3<34> q3<35> q3<36> q3<37> q3<38> q3<39> q3<40> q3<41> 
+ q3<42> q3<43> q3<44> q3<45> q3<46> q3<47> q3<48> q3<49> q3<50> q3<51> q3<52> 
+ q3<53> q3<54> q3<55> q3<56> q3<57> q3<58> q3<59> q3<60> q3<61> q3<62> q3<63> 
+ sl<4> sl<5> sl<6> sl<7> vdd vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> 
+ wl<7> wl<8> wl<9> wl<10> wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> 
+ wl<18> wl<19> wl<20> wl<21> wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> 
+ wl<29> wl<30> wl<31> / inputcell
XI1 bl<0> bl<1> bl<2> bl<3> q0<0> q0<1> q0<2> q0<3> q0<4> q0<5> q0<6> q0<7> 
+ q0<8> q0<9> q0<10> q0<11> q0<12> q0<13> q0<14> q0<15> q0<16> q0<17> q0<18> 
+ q0<19> q0<20> q0<21> q0<22> q0<23> q0<24> q0<25> q0<26> q0<27> q0<28> q0<29> 
+ q0<30> q0<31> q1<0> q1<1> q1<2> q1<3> q1<4> q1<5> q1<6> q1<7> q1<8> q1<9> 
+ q1<10> q1<11> q1<12> q1<13> q1<14> q1<15> q1<16> q1<17> q1<18> q1<19> q1<20> 
+ q1<21> q1<22> q1<23> q1<24> q1<25> q1<26> q1<27> q1<28> q1<29> q1<30> q1<31> 
+ q2<0> q2<1> q2<2> q2<3> q2<4> q2<5> q2<6> q2<7> q2<8> q2<9> q2<10> q2<11> 
+ q2<12> q2<13> q2<14> q2<15> q2<16> q2<17> q2<18> q2<19> q2<20> q2<21> q2<22> 
+ q2<23> q2<24> q2<25> q2<26> q2<27> q2<28> q2<29> q2<30> q2<31> q3<0> q3<1> 
+ q3<2> q3<3> q3<4> q3<5> q3<6> q3<7> q3<8> q3<9> q3<10> q3<11> q3<12> q3<13> 
+ q3<14> q3<15> q3<16> q3<17> q3<18> q3<19> q3<20> q3<21> q3<22> q3<23> q3<24> 
+ q3<25> q3<26> q3<27> q3<28> q3<29> q3<30> q3<31> sl<0> sl<1> sl<2> sl<3> vdd 
+ vss wl<0> wl<1> wl<2> wl<3> wl<4> wl<5> wl<6> wl<7> wl<8> wl<9> wl<10> 
+ wl<11> wl<12> wl<13> wl<14> wl<15> wl<16> wl<17> wl<18> wl<19> wl<20> wl<21> 
+ wl<22> wl<23> wl<24> wl<25> wl<26> wl<27> wl<28> wl<29> wl<30> wl<31> / 
+ inputcell
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    inbuf_decoder
* View Name:    schematic
************************************************************************

.SUBCKT inbuf_decoder a_inbuf<0> a_inbuf<1> a_inbuf<2> a_inbuf<3> a_inbuf<4> 
+ en rowbuf<0> rowbuf<1> rowbuf<2> rowbuf<3> rowbuf<4> rowbuf<5> rowbuf<6> 
+ rowbuf<7> rowbuf<8> rowbuf<9> rowbuf<10> rowbuf<11> rowbuf<12> rowbuf<13> 
+ rowbuf<14> rowbuf<15> rowbuf<16> rowbuf<17> rowbuf<18> rowbuf<19> rowbuf<20> 
+ rowbuf<21> rowbuf<22> rowbuf<23> rowbuf<24> rowbuf<25> rowbuf<26> rowbuf<27> 
+ rowbuf<28> rowbuf<29> rowbuf<30> rowbuf<31> vdd vss
*.PININFO a_inbuf<0>:I a_inbuf<1>:I a_inbuf<2>:I a_inbuf<3>:I a_inbuf<4>:I 
*.PININFO en:I rowbuf<0>:O rowbuf<1>:O rowbuf<2>:O rowbuf<3>:O rowbuf<4>:O 
*.PININFO rowbuf<5>:O rowbuf<6>:O rowbuf<7>:O rowbuf<8>:O rowbuf<9>:O 
*.PININFO rowbuf<10>:O rowbuf<11>:O rowbuf<12>:O rowbuf<13>:O rowbuf<14>:O 
*.PININFO rowbuf<15>:O rowbuf<16>:O rowbuf<17>:O rowbuf<18>:O rowbuf<19>:O 
*.PININFO rowbuf<20>:O rowbuf<21>:O rowbuf<22>:O rowbuf<23>:O rowbuf<24>:O 
*.PININFO rowbuf<25>:O rowbuf<26>:O rowbuf<27>:O rowbuf<28>:O rowbuf<29>:O 
*.PININFO rowbuf<30>:O rowbuf<31>:O vdd:B vss:B
XI6 a_inbuf4b a_inbuf4bn vdd vss / inv1
XI5 net03 a_inbuf4b vdd vss / inv1
XI3 vdd vss a_inbuf4bn a_inbuf<0> a_inbuf<1> a_inbuf<2> a_inbuf<3> rowbuf<16> 
+ rowbuf<17> rowbuf<18> rowbuf<19> rowbuf<20> rowbuf<21> rowbuf<22> rowbuf<23> 
+ rowbuf<24> rowbuf<25> rowbuf<26> rowbuf<27> rowbuf<28> rowbuf<29> rowbuf<30> 
+ rowbuf<31> / 4x16decoder
XI1 vdd vss a_inbuf4b a_inbuf<0> a_inbuf<1> a_inbuf<2> a_inbuf<3> rowbuf<0> 
+ rowbuf<1> rowbuf<2> rowbuf<3> rowbuf<4> rowbuf<5> rowbuf<6> rowbuf<7> 
+ rowbuf<8> rowbuf<9> rowbuf<10> rowbuf<11> rowbuf<12> rowbuf<13> rowbuf<14> 
+ rowbuf<15> / 4x16decoder
XI4 a_inbuf<4> en net03 vdd vss / nor
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv0_3
* View Name:    schematic
************************************************************************

.SUBCKT inv0_3 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    delaycell_editable
* View Name:    schematic
************************************************************************

.SUBCKT delaycell_editable VDD VSS in out
*.PININFO in:I out:O VDD:B VSS:B
XI1<0> x<0> x<1> VDD VSS / inv0_3
XI1<1> x<1> x<2> VDD VSS / inv0_3
XI1<2> x<2> x<3> VDD VSS / inv0_3
XI1<3> x<3> x<4> VDD VSS / inv0_3
XI1<4> x<4> x<5> VDD VSS / inv0_3
XI1<5> x<5> x<6> VDD VSS / inv0_3
XI0 in x<0> VDD VSS / inv0_3
XI2 x<6> out VDD VSS / inv1
XPM3<0> x<1> x<0> x<1> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<1> x<2> x<1> x<2> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<2> x<3> x<2> x<3> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<3> x<4> x<3> x<4> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<4> x<5> x<4> x<5> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM3<5> x<6> x<5> x<6> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM4 out x<6> out VDD p12ll_mis_ckt MR=1 L=80n W=400n
XPM2 x<0> in x<0> VDD p12ll_mis_ckt MR=1 L=80n W=400n
XNM6 out x<6> out VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<0> x<1> x<0> x<1> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<1> x<2> x<1> x<2> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<2> x<3> x<2> x<3> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<3> x<4> x<3> x<4> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<4> x<5> x<4> x<5> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM5<5> x<6> x<5> x<6> VSS n12ll_mis_ckt MR=1 L=80n W=400n
XNM0 x<0> in x<0> VSS n12ll_mis_ckt MR=1 L=80n W=400n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    Tgenerate
* View Name:    schematic
************************************************************************

.SUBCKT Tgenerate en in1 in2 q<0> q<1> q<2> q<3> time<0> time<1> time<2> 
+ time<3> vdd vss
*.PININFO en:I q<0>:I q<1>:I q<2>:I q<3>:I time<0>:I time<1>:I time<2>:I 
*.PININFO time<3>:I in1:O in2:O vdd:B vss:B
XI21 net014 net013 net025 vdd vss / nor
XI17 net15 net14 net19 vdd vss / nor
XI12 net19 en net18 vdd vss / nor
XI22 net024 net026 vdd vss / inv4
XI13 net027 net17 vdd vss / inv4
XI23 net026 in2 vdd vss / inv8
XI14 net17 in1 vdd vss / inv8
XI20 net013 net014 net027 vdd vss / nand
XI7 q<3> time<3> net10 vdd vss / nand
XI6 q<2> time<2> net11 vdd vss / nand
XI16 net11 net10 net14 vdd vss / nand
XI3 q<1> time<1> net12 vdd vss / nand
XI15 net13 net12 net15 vdd vss / nand
XI0 q<0> time<0> net13 vdd vss / nand
XI24 net025 net024 vdd vss / inv1
XI19 net18 net013 vdd vss / inv1
XI27 vdd vss net013 net014 / delaycell_editable
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    timegenerate
* View Name:    schematic
************************************************************************

.SUBCKT timegenerate blbuf<0> blbuf<1> blbuf<2> blbuf<3> blbuf<4> blbuf<5> 
+ blbuf<6> blbuf<7> blbuf<8> blbuf<9> blbuf<10> blbuf<11> blbuf<12> blbuf<13> 
+ blbuf<14> blbuf<15> en in1<0> in1<1> in1<2> in1<3> in1<4> in1<5> in1<6> 
+ in1<7> in1<8> in1<9> in1<10> in1<11> in1<12> in1<13> in1<14> in1<15> in1<16> 
+ in1<17> in1<18> in1<19> in1<20> in1<21> in1<22> in1<23> in1<24> in1<25> 
+ in1<26> in1<27> in1<28> in1<29> in1<30> in1<31> in1<32> in1<33> in1<34> 
+ in1<35> in1<36> in1<37> in1<38> in1<39> in1<40> in1<41> in1<42> in1<43> 
+ in1<44> in1<45> in1<46> in1<47> in1<48> in1<49> in1<50> in1<51> in1<52> 
+ in1<53> in1<54> in1<55> in1<56> in1<57> in1<58> in1<59> in1<60> in1<61> 
+ in1<62> in1<63> in1<64> in1<65> in1<66> in1<67> in1<68> in1<69> in1<70> 
+ in1<71> in1<72> in1<73> in1<74> in1<75> in1<76> in1<77> in1<78> in1<79> 
+ in1<80> in1<81> in1<82> in1<83> in1<84> in1<85> in1<86> in1<87> in1<88> 
+ in1<89> in1<90> in1<91> in1<92> in1<93> in1<94> in1<95> in1<96> in1<97> 
+ in1<98> in1<99> in1<100> in1<101> in1<102> in1<103> in1<104> in1<105> 
+ in1<106> in1<107> in1<108> in1<109> in1<110> in1<111> in1<112> in1<113> 
+ in1<114> in1<115> in1<116> in1<117> in1<118> in1<119> in1<120> in1<121> 
+ in1<122> in1<123> in1<124> in1<125> in1<126> in1<127> in2<0> in2<1> in2<2> 
+ in2<3> in2<4> in2<5> in2<6> in2<7> in2<8> in2<9> in2<10> in2<11> in2<12> 
+ in2<13> in2<14> in2<15> in2<16> in2<17> in2<18> in2<19> in2<20> in2<21> 
+ in2<22> in2<23> in2<24> in2<25> in2<26> in2<27> in2<28> in2<29> in2<30> 
+ in2<31> in2<32> in2<33> in2<34> in2<35> in2<36> in2<37> in2<38> in2<39> 
+ in2<40> in2<41> in2<42> in2<43> in2<44> in2<45> in2<46> in2<47> in2<48> 
+ in2<49> in2<50> in2<51> in2<52> in2<53> in2<54> in2<55> in2<56> in2<57> 
+ in2<58> in2<59> in2<60> in2<61> in2<62> in2<63> in2<64> in2<65> in2<66> 
+ in2<67> in2<68> in2<69> in2<70> in2<71> in2<72> in2<73> in2<74> in2<75> 
+ in2<76> in2<77> in2<78> in2<79> in2<80> in2<81> in2<82> in2<83> in2<84> 
+ in2<85> in2<86> in2<87> in2<88> in2<89> in2<90> in2<91> in2<92> in2<93> 
+ in2<94> in2<95> in2<96> in2<97> in2<98> in2<99> in2<100> in2<101> in2<102> 
+ in2<103> in2<104> in2<105> in2<106> in2<107> in2<108> in2<109> in2<110> 
+ in2<111> in2<112> in2<113> in2<114> in2<115> in2<116> in2<117> in2<118> 
+ in2<119> in2<120> in2<121> in2<122> in2<123> in2<124> in2<125> in2<126> 
+ in2<127> q0<0> q0<1> q0<2> q0<3> q0<4> q0<5> q0<6> q0<7> q0<8> q0<9> q0<10> 
+ q0<11> q0<12> q0<13> q0<14> q0<15> q0<16> q0<17> q0<18> q0<19> q0<20> q0<21> 
+ q0<22> q0<23> q0<24> q0<25> q0<26> q0<27> q0<28> q0<29> q0<30> q0<31> q0<32> 
+ q0<33> q0<34> q0<35> q0<36> q0<37> q0<38> q0<39> q0<40> q0<41> q0<42> q0<43> 
+ q0<44> q0<45> q0<46> q0<47> q0<48> q0<49> q0<50> q0<51> q0<52> q0<53> q0<54> 
+ q0<55> q0<56> q0<57> q0<58> q0<59> q0<60> q0<61> q0<62> q0<63> q0<64> q0<65> 
+ q0<66> q0<67> q0<68> q0<69> q0<70> q0<71> q0<72> q0<73> q0<74> q0<75> q0<76> 
+ q0<77> q0<78> q0<79> q0<80> q0<81> q0<82> q0<83> q0<84> q0<85> q0<86> q0<87> 
+ q0<88> q0<89> q0<90> q0<91> q0<92> q0<93> q0<94> q0<95> q0<96> q0<97> q0<98> 
+ q0<99> q0<100> q0<101> q0<102> q0<103> q0<104> q0<105> q0<106> q0<107> 
+ q0<108> q0<109> q0<110> q0<111> q0<112> q0<113> q0<114> q0<115> q0<116> 
+ q0<117> q0<118> q0<119> q0<120> q0<121> q0<122> q0<123> q0<124> q0<125> 
+ q0<126> q0<127> q1<0> q1<1> q1<2> q1<3> q1<4> q1<5> q1<6> q1<7> q1<8> q1<9> 
+ q1<10> q1<11> q1<12> q1<13> q1<14> q1<15> q1<16> q1<17> q1<18> q1<19> q1<20> 
+ q1<21> q1<22> q1<23> q1<24> q1<25> q1<26> q1<27> q1<28> q1<29> q1<30> q1<31> 
+ q1<32> q1<33> q1<34> q1<35> q1<36> q1<37> q1<38> q1<39> q1<40> q1<41> q1<42> 
+ q1<43> q1<44> q1<45> q1<46> q1<47> q1<48> q1<49> q1<50> q1<51> q1<52> q1<53> 
+ q1<54> q1<55> q1<56> q1<57> q1<58> q1<59> q1<60> q1<61> q1<62> q1<63> q1<64> 
+ q1<65> q1<66> q1<67> q1<68> q1<69> q1<70> q1<71> q1<72> q1<73> q1<74> q1<75> 
+ q1<76> q1<77> q1<78> q1<79> q1<80> q1<81> q1<82> q1<83> q1<84> q1<85> q1<86> 
+ q1<87> q1<88> q1<89> q1<90> q1<91> q1<92> q1<93> q1<94> q1<95> q1<96> q1<97> 
+ q1<98> q1<99> q1<100> q1<101> q1<102> q1<103> q1<104> q1<105> q1<106> 
+ q1<107> q1<108> q1<109> q1<110> q1<111> q1<112> q1<113> q1<114> q1<115> 
+ q1<116> q1<117> q1<118> q1<119> q1<120> q1<121> q1<122> q1<123> q1<124> 
+ q1<125> q1<126> q1<127> q2<0> q2<1> q2<2> q2<3> q2<4> q2<5> q2<6> q2<7> 
+ q2<8> q2<9> q2<10> q2<11> q2<12> q2<13> q2<14> q2<15> q2<16> q2<17> q2<18> 
+ q2<19> q2<20> q2<21> q2<22> q2<23> q2<24> q2<25> q2<26> q2<27> q2<28> q2<29> 
+ q2<30> q2<31> q2<32> q2<33> q2<34> q2<35> q2<36> q2<37> q2<38> q2<39> q2<40> 
+ q2<41> q2<42> q2<43> q2<44> q2<45> q2<46> q2<47> q2<48> q2<49> q2<50> q2<51> 
+ q2<52> q2<53> q2<54> q2<55> q2<56> q2<57> q2<58> q2<59> q2<60> q2<61> q2<62> 
+ q2<63> q2<64> q2<65> q2<66> q2<67> q2<68> q2<69> q2<70> q2<71> q2<72> q2<73> 
+ q2<74> q2<75> q2<76> q2<77> q2<78> q2<79> q2<80> q2<81> q2<82> q2<83> q2<84> 
+ q2<85> q2<86> q2<87> q2<88> q2<89> q2<90> q2<91> q2<92> q2<93> q2<94> q2<95> 
+ q2<96> q2<97> q2<98> q2<99> q2<100> q2<101> q2<102> q2<103> q2<104> q2<105> 
+ q2<106> q2<107> q2<108> q2<109> q2<110> q2<111> q2<112> q2<113> q2<114> 
+ q2<115> q2<116> q2<117> q2<118> q2<119> q2<120> q2<121> q2<122> q2<123> 
+ q2<124> q2<125> q2<126> q2<127> q3<0> q3<1> q3<2> q3<3> q3<4> q3<5> q3<6> 
+ q3<7> q3<8> q3<9> q3<10> q3<11> q3<12> q3<13> q3<14> q3<15> q3<16> q3<17> 
+ q3<18> q3<19> q3<20> q3<21> q3<22> q3<23> q3<24> q3<25> q3<26> q3<27> q3<28> 
+ q3<29> q3<30> q3<31> q3<32> q3<33> q3<34> q3<35> q3<36> q3<37> q3<38> q3<39> 
+ q3<40> q3<41> q3<42> q3<43> q3<44> q3<45> q3<46> q3<47> q3<48> q3<49> q3<50> 
+ q3<51> q3<52> q3<53> q3<54> q3<55> q3<56> q3<57> q3<58> q3<59> q3<60> q3<61> 
+ q3<62> q3<63> q3<64> q3<65> q3<66> q3<67> q3<68> q3<69> q3<70> q3<71> q3<72> 
+ q3<73> q3<74> q3<75> q3<76> q3<77> q3<78> q3<79> q3<80> q3<81> q3<82> q3<83> 
+ q3<84> q3<85> q3<86> q3<87> q3<88> q3<89> q3<90> q3<91> q3<92> q3<93> q3<94> 
+ q3<95> q3<96> q3<97> q3<98> q3<99> q3<100> q3<101> q3<102> q3<103> q3<104> 
+ q3<105> q3<106> q3<107> q3<108> q3<109> q3<110> q3<111> q3<112> q3<113> 
+ q3<114> q3<115> q3<116> q3<117> q3<118> q3<119> q3<120> q3<121> q3<122> 
+ q3<123> q3<124> q3<125> q3<126> q3<127> slbuf<0> slbuf<1> slbuf<2> slbuf<3> 
+ slbuf<4> slbuf<5> slbuf<6> slbuf<7> slbuf<8> slbuf<9> slbuf<10> slbuf<11> 
+ slbuf<12> slbuf<13> slbuf<14> slbuf<15> time<0> time<1> time<2> time<3> vdd 
+ vss
*.PININFO en:I q0<0>:I q0<1>:I q0<2>:I q0<3>:I q0<4>:I q0<5>:I q0<6>:I q0<7>:I 
*.PININFO q0<8>:I q0<9>:I q0<10>:I q0<11>:I q0<12>:I q0<13>:I q0<14>:I 
*.PININFO q0<15>:I q0<16>:I q0<17>:I q0<18>:I q0<19>:I q0<20>:I q0<21>:I 
*.PININFO q0<22>:I q0<23>:I q0<24>:I q0<25>:I q0<26>:I q0<27>:I q0<28>:I 
*.PININFO q0<29>:I q0<30>:I q0<31>:I q0<32>:I q0<33>:I q0<34>:I q0<35>:I 
*.PININFO q0<36>:I q0<37>:I q0<38>:I q0<39>:I q0<40>:I q0<41>:I q0<42>:I 
*.PININFO q0<43>:I q0<44>:I q0<45>:I q0<46>:I q0<47>:I q0<48>:I q0<49>:I 
*.PININFO q0<50>:I q0<51>:I q0<52>:I q0<53>:I q0<54>:I q0<55>:I q0<56>:I 
*.PININFO q0<57>:I q0<58>:I q0<59>:I q0<60>:I q0<61>:I q0<62>:I q0<63>:I 
*.PININFO q0<64>:I q0<65>:I q0<66>:I q0<67>:I q0<68>:I q0<69>:I q0<70>:I 
*.PININFO q0<71>:I q0<72>:I q0<73>:I q0<74>:I q0<75>:I q0<76>:I q0<77>:I 
*.PININFO q0<78>:I q0<79>:I q0<80>:I q0<81>:I q0<82>:I q0<83>:I q0<84>:I 
*.PININFO q0<85>:I q0<86>:I q0<87>:I q0<88>:I q0<89>:I q0<90>:I q0<91>:I 
*.PININFO q0<92>:I q0<93>:I q0<94>:I q0<95>:I q0<96>:I q0<97>:I q0<98>:I 
*.PININFO q0<99>:I q0<100>:I q0<101>:I q0<102>:I q0<103>:I q0<104>:I q0<105>:I 
*.PININFO q0<106>:I q0<107>:I q0<108>:I q0<109>:I q0<110>:I q0<111>:I 
*.PININFO q0<112>:I q0<113>:I q0<114>:I q0<115>:I q0<116>:I q0<117>:I 
*.PININFO q0<118>:I q0<119>:I q0<120>:I q0<121>:I q0<122>:I q0<123>:I 
*.PININFO q0<124>:I q0<125>:I q0<126>:I q0<127>:I q1<0>:I q1<1>:I q1<2>:I 
*.PININFO q1<3>:I q1<4>:I q1<5>:I q1<6>:I q1<7>:I q1<8>:I q1<9>:I q1<10>:I 
*.PININFO q1<11>:I q1<12>:I q1<13>:I q1<14>:I q1<15>:I q1<16>:I q1<17>:I 
*.PININFO q1<18>:I q1<19>:I q1<20>:I q1<21>:I q1<22>:I q1<23>:I q1<24>:I 
*.PININFO q1<25>:I q1<26>:I q1<27>:I q1<28>:I q1<29>:I q1<30>:I q1<31>:I 
*.PININFO q1<32>:I q1<33>:I q1<34>:I q1<35>:I q1<36>:I q1<37>:I q1<38>:I 
*.PININFO q1<39>:I q1<40>:I q1<41>:I q1<42>:I q1<43>:I q1<44>:I q1<45>:I 
*.PININFO q1<46>:I q1<47>:I q1<48>:I q1<49>:I q1<50>:I q1<51>:I q1<52>:I 
*.PININFO q1<53>:I q1<54>:I q1<55>:I q1<56>:I q1<57>:I q1<58>:I q1<59>:I 
*.PININFO q1<60>:I q1<61>:I q1<62>:I q1<63>:I q1<64>:I q1<65>:I q1<66>:I 
*.PININFO q1<67>:I q1<68>:I q1<69>:I q1<70>:I q1<71>:I q1<72>:I q1<73>:I 
*.PININFO q1<74>:I q1<75>:I q1<76>:I q1<77>:I q1<78>:I q1<79>:I q1<80>:I 
*.PININFO q1<81>:I q1<82>:I q1<83>:I q1<84>:I q1<85>:I q1<86>:I q1<87>:I 
*.PININFO q1<88>:I q1<89>:I q1<90>:I q1<91>:I q1<92>:I q1<93>:I q1<94>:I 
*.PININFO q1<95>:I q1<96>:I q1<97>:I q1<98>:I q1<99>:I q1<100>:I q1<101>:I 
*.PININFO q1<102>:I q1<103>:I q1<104>:I q1<105>:I q1<106>:I q1<107>:I 
*.PININFO q1<108>:I q1<109>:I q1<110>:I q1<111>:I q1<112>:I q1<113>:I 
*.PININFO q1<114>:I q1<115>:I q1<116>:I q1<117>:I q1<118>:I q1<119>:I 
*.PININFO q1<120>:I q1<121>:I q1<122>:I q1<123>:I q1<124>:I q1<125>:I 
*.PININFO q1<126>:I q1<127>:I q2<0>:I q2<1>:I q2<2>:I q2<3>:I q2<4>:I q2<5>:I 
*.PININFO q2<6>:I q2<7>:I q2<8>:I q2<9>:I q2<10>:I q2<11>:I q2<12>:I q2<13>:I 
*.PININFO q2<14>:I q2<15>:I q2<16>:I q2<17>:I q2<18>:I q2<19>:I q2<20>:I 
*.PININFO q2<21>:I q2<22>:I q2<23>:I q2<24>:I q2<25>:I q2<26>:I q2<27>:I 
*.PININFO q2<28>:I q2<29>:I q2<30>:I q2<31>:I q2<32>:I q2<33>:I q2<34>:I 
*.PININFO q2<35>:I q2<36>:I q2<37>:I q2<38>:I q2<39>:I q2<40>:I q2<41>:I 
*.PININFO q2<42>:I q2<43>:I q2<44>:I q2<45>:I q2<46>:I q2<47>:I q2<48>:I 
*.PININFO q2<49>:I q2<50>:I q2<51>:I q2<52>:I q2<53>:I q2<54>:I q2<55>:I 
*.PININFO q2<56>:I q2<57>:I q2<58>:I q2<59>:I q2<60>:I q2<61>:I q2<62>:I 
*.PININFO q2<63>:I q2<64>:I q2<65>:I q2<66>:I q2<67>:I q2<68>:I q2<69>:I 
*.PININFO q2<70>:I q2<71>:I q2<72>:I q2<73>:I q2<74>:I q2<75>:I q2<76>:I 
*.PININFO q2<77>:I q2<78>:I q2<79>:I q2<80>:I q2<81>:I q2<82>:I q2<83>:I 
*.PININFO q2<84>:I q2<85>:I q2<86>:I q2<87>:I q2<88>:I q2<89>:I q2<90>:I 
*.PININFO q2<91>:I q2<92>:I q2<93>:I q2<94>:I q2<95>:I q2<96>:I q2<97>:I 
*.PININFO q2<98>:I q2<99>:I q2<100>:I q2<101>:I q2<102>:I q2<103>:I q2<104>:I 
*.PININFO q2<105>:I q2<106>:I q2<107>:I q2<108>:I q2<109>:I q2<110>:I 
*.PININFO q2<111>:I q2<112>:I q2<113>:I q2<114>:I q2<115>:I q2<116>:I 
*.PININFO q2<117>:I q2<118>:I q2<119>:I q2<120>:I q2<121>:I q2<122>:I 
*.PININFO q2<123>:I q2<124>:I q2<125>:I q2<126>:I q2<127>:I q3<0>:I q3<1>:I 
*.PININFO q3<2>:I q3<3>:I q3<4>:I q3<5>:I q3<6>:I q3<7>:I q3<8>:I q3<9>:I 
*.PININFO q3<10>:I q3<11>:I q3<12>:I q3<13>:I q3<14>:I q3<15>:I q3<16>:I 
*.PININFO q3<17>:I q3<18>:I q3<19>:I q3<20>:I q3<21>:I q3<22>:I q3<23>:I 
*.PININFO q3<24>:I q3<25>:I q3<26>:I q3<27>:I q3<28>:I q3<29>:I q3<30>:I 
*.PININFO q3<31>:I q3<32>:I q3<33>:I q3<34>:I q3<35>:I q3<36>:I q3<37>:I 
*.PININFO q3<38>:I q3<39>:I q3<40>:I q3<41>:I q3<42>:I q3<43>:I q3<44>:I 
*.PININFO q3<45>:I q3<46>:I q3<47>:I q3<48>:I q3<49>:I q3<50>:I q3<51>:I 
*.PININFO q3<52>:I q3<53>:I q3<54>:I q3<55>:I q3<56>:I q3<57>:I q3<58>:I 
*.PININFO q3<59>:I q3<60>:I q3<61>:I q3<62>:I q3<63>:I q3<64>:I q3<65>:I 
*.PININFO q3<66>:I q3<67>:I q3<68>:I q3<69>:I q3<70>:I q3<71>:I q3<72>:I 
*.PININFO q3<73>:I q3<74>:I q3<75>:I q3<76>:I q3<77>:I q3<78>:I q3<79>:I 
*.PININFO q3<80>:I q3<81>:I q3<82>:I q3<83>:I q3<84>:I q3<85>:I q3<86>:I 
*.PININFO q3<87>:I q3<88>:I q3<89>:I q3<90>:I q3<91>:I q3<92>:I q3<93>:I 
*.PININFO q3<94>:I q3<95>:I q3<96>:I q3<97>:I q3<98>:I q3<99>:I q3<100>:I 
*.PININFO q3<101>:I q3<102>:I q3<103>:I q3<104>:I q3<105>:I q3<106>:I 
*.PININFO q3<107>:I q3<108>:I q3<109>:I q3<110>:I q3<111>:I q3<112>:I 
*.PININFO q3<113>:I q3<114>:I q3<115>:I q3<116>:I q3<117>:I q3<118>:I 
*.PININFO q3<119>:I q3<120>:I q3<121>:I q3<122>:I q3<123>:I q3<124>:I 
*.PININFO q3<125>:I q3<126>:I q3<127>:I time<0>:I time<1>:I time<2>:I 
*.PININFO time<3>:I in1<0>:O in1<1>:O in1<2>:O in1<3>:O in1<4>:O in1<5>:O 
*.PININFO in1<6>:O in1<7>:O in1<8>:O in1<9>:O in1<10>:O in1<11>:O in1<12>:O 
*.PININFO in1<13>:O in1<14>:O in1<15>:O in1<16>:O in1<17>:O in1<18>:O 
*.PININFO in1<19>:O in1<20>:O in1<21>:O in1<22>:O in1<23>:O in1<24>:O 
*.PININFO in1<25>:O in1<26>:O in1<27>:O in1<28>:O in1<29>:O in1<30>:O 
*.PININFO in1<31>:O in1<32>:O in1<33>:O in1<34>:O in1<35>:O in1<36>:O 
*.PININFO in1<37>:O in1<38>:O in1<39>:O in1<40>:O in1<41>:O in1<42>:O 
*.PININFO in1<43>:O in1<44>:O in1<45>:O in1<46>:O in1<47>:O in1<48>:O 
*.PININFO in1<49>:O in1<50>:O in1<51>:O in1<52>:O in1<53>:O in1<54>:O 
*.PININFO in1<55>:O in1<56>:O in1<57>:O in1<58>:O in1<59>:O in1<60>:O 
*.PININFO in1<61>:O in1<62>:O in1<63>:O in1<64>:O in1<65>:O in1<66>:O 
*.PININFO in1<67>:O in1<68>:O in1<69>:O in1<70>:O in1<71>:O in1<72>:O 
*.PININFO in1<73>:O in1<74>:O in1<75>:O in1<76>:O in1<77>:O in1<78>:O 
*.PININFO in1<79>:O in1<80>:O in1<81>:O in1<82>:O in1<83>:O in1<84>:O 
*.PININFO in1<85>:O in1<86>:O in1<87>:O in1<88>:O in1<89>:O in1<90>:O 
*.PININFO in1<91>:O in1<92>:O in1<93>:O in1<94>:O in1<95>:O in1<96>:O 
*.PININFO in1<97>:O in1<98>:O in1<99>:O in1<100>:O in1<101>:O in1<102>:O 
*.PININFO in1<103>:O in1<104>:O in1<105>:O in1<106>:O in1<107>:O in1<108>:O 
*.PININFO in1<109>:O in1<110>:O in1<111>:O in1<112>:O in1<113>:O in1<114>:O 
*.PININFO in1<115>:O in1<116>:O in1<117>:O in1<118>:O in1<119>:O in1<120>:O 
*.PININFO in1<121>:O in1<122>:O in1<123>:O in1<124>:O in1<125>:O in1<126>:O 
*.PININFO in1<127>:O in2<0>:O in2<1>:O in2<2>:O in2<3>:O in2<4>:O in2<5>:O 
*.PININFO in2<6>:O in2<7>:O in2<8>:O in2<9>:O in2<10>:O in2<11>:O in2<12>:O 
*.PININFO in2<13>:O in2<14>:O in2<15>:O in2<16>:O in2<17>:O in2<18>:O 
*.PININFO in2<19>:O in2<20>:O in2<21>:O in2<22>:O in2<23>:O in2<24>:O 
*.PININFO in2<25>:O in2<26>:O in2<27>:O in2<28>:O in2<29>:O in2<30>:O 
*.PININFO in2<31>:O in2<32>:O in2<33>:O in2<34>:O in2<35>:O in2<36>:O 
*.PININFO in2<37>:O in2<38>:O in2<39>:O in2<40>:O in2<41>:O in2<42>:O 
*.PININFO in2<43>:O in2<44>:O in2<45>:O in2<46>:O in2<47>:O in2<48>:O 
*.PININFO in2<49>:O in2<50>:O in2<51>:O in2<52>:O in2<53>:O in2<54>:O 
*.PININFO in2<55>:O in2<56>:O in2<57>:O in2<58>:O in2<59>:O in2<60>:O 
*.PININFO in2<61>:O in2<62>:O in2<63>:O in2<64>:O in2<65>:O in2<66>:O 
*.PININFO in2<67>:O in2<68>:O in2<69>:O in2<70>:O in2<71>:O in2<72>:O 
*.PININFO in2<73>:O in2<74>:O in2<75>:O in2<76>:O in2<77>:O in2<78>:O 
*.PININFO in2<79>:O in2<80>:O in2<81>:O in2<82>:O in2<83>:O in2<84>:O 
*.PININFO in2<85>:O in2<86>:O in2<87>:O in2<88>:O in2<89>:O in2<90>:O 
*.PININFO in2<91>:O in2<92>:O in2<93>:O in2<94>:O in2<95>:O in2<96>:O 
*.PININFO in2<97>:O in2<98>:O in2<99>:O in2<100>:O in2<101>:O in2<102>:O 
*.PININFO in2<103>:O in2<104>:O in2<105>:O in2<106>:O in2<107>:O in2<108>:O 
*.PININFO in2<109>:O in2<110>:O in2<111>:O in2<112>:O in2<113>:O in2<114>:O 
*.PININFO in2<115>:O in2<116>:O in2<117>:O in2<118>:O in2<119>:O in2<120>:O 
*.PININFO in2<121>:O in2<122>:O in2<123>:O in2<124>:O in2<125>:O in2<126>:O 
*.PININFO in2<127>:O blbuf<0>:B blbuf<1>:B blbuf<2>:B blbuf<3>:B blbuf<4>:B 
*.PININFO blbuf<5>:B blbuf<6>:B blbuf<7>:B blbuf<8>:B blbuf<9>:B blbuf<10>:B 
*.PININFO blbuf<11>:B blbuf<12>:B blbuf<13>:B blbuf<14>:B blbuf<15>:B 
*.PININFO slbuf<0>:B slbuf<1>:B slbuf<2>:B slbuf<3>:B slbuf<4>:B slbuf<5>:B 
*.PININFO slbuf<6>:B slbuf<7>:B slbuf<8>:B slbuf<9>:B slbuf<10>:B slbuf<11>:B 
*.PININFO slbuf<12>:B slbuf<13>:B slbuf<14>:B slbuf<15>:B vdd:B vss:B
XI0<0> enb in1<0> in2<0> q0<0> q1<0> q2<0> q3<0> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<1> enb in1<1> in2<1> q0<1> q1<1> q2<1> q3<1> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<2> enb in1<2> in2<2> q0<2> q1<2> q2<2> q3<2> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<3> enb in1<3> in2<3> q0<3> q1<3> q2<3> q3<3> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<4> enb in1<4> in2<4> q0<4> q1<4> q2<4> q3<4> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<5> enb in1<5> in2<5> q0<5> q1<5> q2<5> q3<5> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<6> enb in1<6> in2<6> q0<6> q1<6> q2<6> q3<6> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<7> enb in1<7> in2<7> q0<7> q1<7> q2<7> q3<7> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<8> enb in1<8> in2<8> q0<8> q1<8> q2<8> q3<8> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<9> enb in1<9> in2<9> q0<9> q1<9> q2<9> q3<9> timeb<0> timeb<1> timeb<2> 
+ timeb<3> vdd vss / Tgenerate
XI0<10> enb in1<10> in2<10> q0<10> q1<10> q2<10> q3<10> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<11> enb in1<11> in2<11> q0<11> q1<11> q2<11> q3<11> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<12> enb in1<12> in2<12> q0<12> q1<12> q2<12> q3<12> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<13> enb in1<13> in2<13> q0<13> q1<13> q2<13> q3<13> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<14> enb in1<14> in2<14> q0<14> q1<14> q2<14> q3<14> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<15> enb in1<15> in2<15> q0<15> q1<15> q2<15> q3<15> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<16> enb in1<16> in2<16> q0<16> q1<16> q2<16> q3<16> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<17> enb in1<17> in2<17> q0<17> q1<17> q2<17> q3<17> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<18> enb in1<18> in2<18> q0<18> q1<18> q2<18> q3<18> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<19> enb in1<19> in2<19> q0<19> q1<19> q2<19> q3<19> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<20> enb in1<20> in2<20> q0<20> q1<20> q2<20> q3<20> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<21> enb in1<21> in2<21> q0<21> q1<21> q2<21> q3<21> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<22> enb in1<22> in2<22> q0<22> q1<22> q2<22> q3<22> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<23> enb in1<23> in2<23> q0<23> q1<23> q2<23> q3<23> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<24> enb in1<24> in2<24> q0<24> q1<24> q2<24> q3<24> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<25> enb in1<25> in2<25> q0<25> q1<25> q2<25> q3<25> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<26> enb in1<26> in2<26> q0<26> q1<26> q2<26> q3<26> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<27> enb in1<27> in2<27> q0<27> q1<27> q2<27> q3<27> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<28> enb in1<28> in2<28> q0<28> q1<28> q2<28> q3<28> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<29> enb in1<29> in2<29> q0<29> q1<29> q2<29> q3<29> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<30> enb in1<30> in2<30> q0<30> q1<30> q2<30> q3<30> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<31> enb in1<31> in2<31> q0<31> q1<31> q2<31> q3<31> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<32> enb in1<32> in2<32> q0<32> q1<32> q2<32> q3<32> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<33> enb in1<33> in2<33> q0<33> q1<33> q2<33> q3<33> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<34> enb in1<34> in2<34> q0<34> q1<34> q2<34> q3<34> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<35> enb in1<35> in2<35> q0<35> q1<35> q2<35> q3<35> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<36> enb in1<36> in2<36> q0<36> q1<36> q2<36> q3<36> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<37> enb in1<37> in2<37> q0<37> q1<37> q2<37> q3<37> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<38> enb in1<38> in2<38> q0<38> q1<38> q2<38> q3<38> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<39> enb in1<39> in2<39> q0<39> q1<39> q2<39> q3<39> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<40> enb in1<40> in2<40> q0<40> q1<40> q2<40> q3<40> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<41> enb in1<41> in2<41> q0<41> q1<41> q2<41> q3<41> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<42> enb in1<42> in2<42> q0<42> q1<42> q2<42> q3<42> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<43> enb in1<43> in2<43> q0<43> q1<43> q2<43> q3<43> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<44> enb in1<44> in2<44> q0<44> q1<44> q2<44> q3<44> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<45> enb in1<45> in2<45> q0<45> q1<45> q2<45> q3<45> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<46> enb in1<46> in2<46> q0<46> q1<46> q2<46> q3<46> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<47> enb in1<47> in2<47> q0<47> q1<47> q2<47> q3<47> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<48> enb in1<48> in2<48> q0<48> q1<48> q2<48> q3<48> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<49> enb in1<49> in2<49> q0<49> q1<49> q2<49> q3<49> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<50> enb in1<50> in2<50> q0<50> q1<50> q2<50> q3<50> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<51> enb in1<51> in2<51> q0<51> q1<51> q2<51> q3<51> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<52> enb in1<52> in2<52> q0<52> q1<52> q2<52> q3<52> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<53> enb in1<53> in2<53> q0<53> q1<53> q2<53> q3<53> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<54> enb in1<54> in2<54> q0<54> q1<54> q2<54> q3<54> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<55> enb in1<55> in2<55> q0<55> q1<55> q2<55> q3<55> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<56> enb in1<56> in2<56> q0<56> q1<56> q2<56> q3<56> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<57> enb in1<57> in2<57> q0<57> q1<57> q2<57> q3<57> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<58> enb in1<58> in2<58> q0<58> q1<58> q2<58> q3<58> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<59> enb in1<59> in2<59> q0<59> q1<59> q2<59> q3<59> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<60> enb in1<60> in2<60> q0<60> q1<60> q2<60> q3<60> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<61> enb in1<61> in2<61> q0<61> q1<61> q2<61> q3<61> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<62> enb in1<62> in2<62> q0<62> q1<62> q2<62> q3<62> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<63> enb in1<63> in2<63> q0<63> q1<63> q2<63> q3<63> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<64> enb in1<64> in2<64> q0<64> q1<64> q2<64> q3<64> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<65> enb in1<65> in2<65> q0<65> q1<65> q2<65> q3<65> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<66> enb in1<66> in2<66> q0<66> q1<66> q2<66> q3<66> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<67> enb in1<67> in2<67> q0<67> q1<67> q2<67> q3<67> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<68> enb in1<68> in2<68> q0<68> q1<68> q2<68> q3<68> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<69> enb in1<69> in2<69> q0<69> q1<69> q2<69> q3<69> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<70> enb in1<70> in2<70> q0<70> q1<70> q2<70> q3<70> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<71> enb in1<71> in2<71> q0<71> q1<71> q2<71> q3<71> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<72> enb in1<72> in2<72> q0<72> q1<72> q2<72> q3<72> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<73> enb in1<73> in2<73> q0<73> q1<73> q2<73> q3<73> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<74> enb in1<74> in2<74> q0<74> q1<74> q2<74> q3<74> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<75> enb in1<75> in2<75> q0<75> q1<75> q2<75> q3<75> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<76> enb in1<76> in2<76> q0<76> q1<76> q2<76> q3<76> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<77> enb in1<77> in2<77> q0<77> q1<77> q2<77> q3<77> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<78> enb in1<78> in2<78> q0<78> q1<78> q2<78> q3<78> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<79> enb in1<79> in2<79> q0<79> q1<79> q2<79> q3<79> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<80> enb in1<80> in2<80> q0<80> q1<80> q2<80> q3<80> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<81> enb in1<81> in2<81> q0<81> q1<81> q2<81> q3<81> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<82> enb in1<82> in2<82> q0<82> q1<82> q2<82> q3<82> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<83> enb in1<83> in2<83> q0<83> q1<83> q2<83> q3<83> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<84> enb in1<84> in2<84> q0<84> q1<84> q2<84> q3<84> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<85> enb in1<85> in2<85> q0<85> q1<85> q2<85> q3<85> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<86> enb in1<86> in2<86> q0<86> q1<86> q2<86> q3<86> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<87> enb in1<87> in2<87> q0<87> q1<87> q2<87> q3<87> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<88> enb in1<88> in2<88> q0<88> q1<88> q2<88> q3<88> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<89> enb in1<89> in2<89> q0<89> q1<89> q2<89> q3<89> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<90> enb in1<90> in2<90> q0<90> q1<90> q2<90> q3<90> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<91> enb in1<91> in2<91> q0<91> q1<91> q2<91> q3<91> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<92> enb in1<92> in2<92> q0<92> q1<92> q2<92> q3<92> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<93> enb in1<93> in2<93> q0<93> q1<93> q2<93> q3<93> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<94> enb in1<94> in2<94> q0<94> q1<94> q2<94> q3<94> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<95> enb in1<95> in2<95> q0<95> q1<95> q2<95> q3<95> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<96> enb in1<96> in2<96> q0<96> q1<96> q2<96> q3<96> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<97> enb in1<97> in2<97> q0<97> q1<97> q2<97> q3<97> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<98> enb in1<98> in2<98> q0<98> q1<98> q2<98> q3<98> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<99> enb in1<99> in2<99> q0<99> q1<99> q2<99> q3<99> timeb<0> timeb<1> 
+ timeb<2> timeb<3> vdd vss / Tgenerate
XI0<100> enb in1<100> in2<100> q0<100> q1<100> q2<100> q3<100> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<101> enb in1<101> in2<101> q0<101> q1<101> q2<101> q3<101> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<102> enb in1<102> in2<102> q0<102> q1<102> q2<102> q3<102> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<103> enb in1<103> in2<103> q0<103> q1<103> q2<103> q3<103> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<104> enb in1<104> in2<104> q0<104> q1<104> q2<104> q3<104> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<105> enb in1<105> in2<105> q0<105> q1<105> q2<105> q3<105> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<106> enb in1<106> in2<106> q0<106> q1<106> q2<106> q3<106> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<107> enb in1<107> in2<107> q0<107> q1<107> q2<107> q3<107> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<108> enb in1<108> in2<108> q0<108> q1<108> q2<108> q3<108> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<109> enb in1<109> in2<109> q0<109> q1<109> q2<109> q3<109> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<110> enb in1<110> in2<110> q0<110> q1<110> q2<110> q3<110> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<111> enb in1<111> in2<111> q0<111> q1<111> q2<111> q3<111> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<112> enb in1<112> in2<112> q0<112> q1<112> q2<112> q3<112> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<113> enb in1<113> in2<113> q0<113> q1<113> q2<113> q3<113> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<114> enb in1<114> in2<114> q0<114> q1<114> q2<114> q3<114> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<115> enb in1<115> in2<115> q0<115> q1<115> q2<115> q3<115> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<116> enb in1<116> in2<116> q0<116> q1<116> q2<116> q3<116> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<117> enb in1<117> in2<117> q0<117> q1<117> q2<117> q3<117> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<118> enb in1<118> in2<118> q0<118> q1<118> q2<118> q3<118> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<119> enb in1<119> in2<119> q0<119> q1<119> q2<119> q3<119> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<120> enb in1<120> in2<120> q0<120> q1<120> q2<120> q3<120> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<121> enb in1<121> in2<121> q0<121> q1<121> q2<121> q3<121> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<122> enb in1<122> in2<122> q0<122> q1<122> q2<122> q3<122> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<123> enb in1<123> in2<123> q0<123> q1<123> q2<123> q3<123> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<124> enb in1<124> in2<124> q0<124> q1<124> q2<124> q3<124> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<125> enb in1<125> in2<125> q0<125> q1<125> q2<125> q3<125> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<126> enb in1<126> in2<126> q0<126> q1<126> q2<126> q3<126> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI0<127> enb in1<127> in2<127> q0<127> q1<127> q2<127> q3<127> timeb<0> 
+ timeb<1> timeb<2> timeb<3> vdd vss / Tgenerate
XI2 net09 enb vdd vss / inv8
XI1<0> net019<0> timeb<0> vdd vss / inv8
XI1<1> net019<1> timeb<1> vdd vss / inv8
XI1<2> net019<2> timeb<2> vdd vss / inv8
XI1<3> net019<3> timeb<3> vdd vss / inv8
XI3 en net09 vdd vss / inv4
XI25<0> time<0> net019<0> vdd vss / inv4
XI25<1> time<1> net019<1> vdd vss / inv4
XI25<2> time<2> net019<2> vdd vss / inv4
XI25<3> time<3> net019<3> vdd vss / inv4
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    Dtriger
* View Name:    schematic
************************************************************************

.SUBCKT Dtriger cp d q qn rdn sdn vdd vss
*.PININFO cp:I d:I rdn:I sdn:I q:O qn:O vdd:B vss:B
XI12 vdd vss net10 sdn net19 net27 / 3nand
XI9 vdd vss rdn net27 cp net19 / 3nand
XI8 vdd vss qn net19 sdn q / 3nand
XI11 vdd vss net18 rdn d net10 / 3nand
XI6 vdd vss rdn net18 q qn / 3nand
XI10 vdd vss cp net10 net19 net18 / 3nand
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    countercell
* View Name:    schematic
************************************************************************

.SUBCKT countercell cp q<0> q<1> q<2> q<3> q<4> q<5> setn vdd vss
*.PININFO cp:I setn:I q<0>:O q<1>:O q<2>:O q<3>:O q<4>:O q<5>:O vdd:B vss:B
XI14 net67 net69 net70 net69 setn vdd vdd vss / Dtriger
XI13 net65 net67 net68 net67 setn vdd vdd vss / Dtriger
XI12 net61 net63 net64 net63 setn vdd vdd vss / Dtriger
XI11 net63 net65 net66 net65 setn vdd vdd vss / Dtriger
XI8 net59 net61 net62 net61 setn vdd vdd vss / Dtriger
XI0 cp net59 net60 net59 setn vdd vdd vss / Dtriger
XI22 net72 q<4> vdd vss / inv1
XI21 net73 q<5> vdd vss / inv1
XI20 net74 q<3> vdd vss / inv1
XI19 net75 q<2> vdd vss / inv1
XI18 net76 q<1> vdd vss / inv1
XI17 net77 q<0> vdd vss / inv1
XI16 net68 net72 vdd vss / inv1
XI15 net70 net73 vdd vss / inv1
XI10 net66 net74 vdd vss / inv1
XI9 net64 net75 vdd vss / inv1
XI3 net60 net77 vdd vss / inv1
XI7 net62 net76 vdd vss / inv1
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    inv0_5
* View Name:    schematic
************************************************************************

.SUBCKT inv0_5 IN OUT VDD VSS
*.PININFO IN:B OUT:B VDD:B VSS:B
XPM1 OUT IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XNM1 OUT IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    countercell2
* View Name:    schematic
************************************************************************

.SUBCKT countercell2 adco<0> adco<1> op<0> op<1> op<2> op<3> op<4> op<5> op<6> 
+ op<7> op<8> op<9> op<10> op<11> out setn vdd vss
*.PININFO adco<0>:I adco<1>:I op<0>:I op<1>:I op<2>:I op<3>:I op<4>:I op<5>:I 
*.PININFO op<6>:I op<7>:I op<8>:I op<9>:I op<10>:I op<11>:I setn:I out:O vdd:B 
*.PININFO vss:B
XI1 adco<1> q<6> q<7> q<8> q<9> q<10> q<11> setn vdd vss / countercell
XI0 adco<0> q<0> q<1> q<2> q<3> q<4> q<5> setn vdd vss / countercell
XI2<0> q<0> op<0> net10<0> out vdd vss / Tgate
XI2<1> q<1> op<1> net10<1> out vdd vss / Tgate
XI2<2> q<2> op<2> net10<2> out vdd vss / Tgate
XI2<3> q<3> op<3> net10<3> out vdd vss / Tgate
XI2<4> q<4> op<4> net10<4> out vdd vss / Tgate
XI2<5> q<5> op<5> net10<5> out vdd vss / Tgate
XI2<6> q<6> op<6> net10<6> out vdd vss / Tgate
XI2<7> q<7> op<7> net10<7> out vdd vss / Tgate
XI2<8> q<8> op<8> net10<8> out vdd vss / Tgate
XI2<9> q<9> op<9> net10<9> out vdd vss / Tgate
XI2<10> q<10> op<10> net10<10> out vdd vss / Tgate
XI2<11> q<11> op<11> net10<11> out vdd vss / Tgate
XI3<0> op<0> net10<0> vdd vss / inv0_5
XI3<1> op<1> net10<1> vdd vss / inv0_5
XI3<2> op<2> net10<2> vdd vss / inv0_5
XI3<3> op<3> net10<3> vdd vss / inv0_5
XI3<4> op<4> net10<4> vdd vss / inv0_5
XI3<5> op<5> net10<5> vdd vss / inv0_5
XI3<6> op<6> net10<6> vdd vss / inv0_5
XI3<7> op<7> net10<7> vdd vss / inv0_5
XI3<8> op<8> net10<8> vdd vss / inv0_5
XI3<9> op<9> net10<9> vdd vss / inv0_5
XI3<10> op<10> net10<10> vdd vss / inv0_5
XI3<11> op<11> net10<11> vdd vss / inv0_5
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    4x16decoder2
* View Name:    schematic
************************************************************************

.SUBCKT 4x16decoder2 VDD VSS en in<0> in<1> in<2> in<3> out<0> out<1> out<2> 
+ out<3> out<4> out<5> out<6> out<7> out<8> out<9> out<10> out<11> out<12> 
+ out<13> out<14> out<15>
*.PININFO en:I in<0>:I in<1>:I in<2>:I in<3>:I out<0>:O out<1>:O out<2>:O 
*.PININFO out<3>:O out<4>:O out<5>:O out<6>:O out<7>:O out<8>:O out<9>:O 
*.PININFO out<10>:O out<11>:O out<12>:O out<13>:O out<14>:O out<15>:O VDD:B 
*.PININFO VSS:B
XI15 VDD VSS en in<2> in<3> b<0> b<1> b<2> b<3> / 2x4decoder
XI0 VDD VSS en in<0> in<1> c<0> c<1> c<2> c<3> / 2x4decoder
XI73 net173 out<15> VDD VSS / inv4
XI70 net174 out<14> VDD VSS / inv4
XI69 net175 out<13> VDD VSS / inv4
XI67 net176 out<12> VDD VSS / inv4
XI81 net092 out<11> VDD VSS / inv4
XI78 net097 out<10> VDD VSS / inv4
XI77 net179 out<9> VDD VSS / inv4
XI75 net180 out<8> VDD VSS / inv4
XI65 net0112 out<7> VDD VSS / inv4
XI62 net182 out<6> VDD VSS / inv4
XI61 net183 out<5> VDD VSS / inv4
XI59 net0127 out<4> VDD VSS / inv4
XI57 net185 out<3> VDD VSS / inv4
XI54 net0137 out<2> VDD VSS / inv4
XI53 net187 out<1> VDD VSS / inv4
XI51 net188 out<0> VDD VSS / inv4
XI8 c<2> b<2> net097 VDD VSS / nand
XI7 c<3> b<2> net092 VDD VSS / nand
XI6 c<3> b<1> net0112 VDD VSS / nand
XI5 c<2> b<1> net182 VDD VSS / nand
XI4 c<0> b<1> net0127 VDD VSS / nand
XI3 c<1> b<1> net183 VDD VSS / nand
XI2 c<3> b<0> net185 VDD VSS / nand
XI1 c<2> b<0> net0137 VDD VSS / nand
XI9 c<0> b<2> net180 VDD VSS / nand
XI10 c<1> b<2> net179 VDD VSS / nand
XI11 c<1> b<3> net175 VDD VSS / nand
XI12 c<0> b<3> net176 VDD VSS / nand
XI13 c<2> b<3> net174 VDD VSS / nand
XI14 c<3> b<3> net173 VDD VSS / nand
XI50 c<0> b<0> net188 VDD VSS / nand
XI52 c<1> b<0> net187 VDD VSS / nand
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    counter
* View Name:    schematic
************************************************************************

.SUBCKT counter a_read<0> a_read<1> a_read<2> a_read<3> adc<0> adc<1> adc<2> 
+ adc<3> adc<4> adc<5> adc<6> adc<7> adc<8> adc<9> adc<10> adc<11> adc<12> 
+ adc<13> adc<14> adc<15> adc<16> adc<17> adc<18> adc<19> adc<20> adc<21> 
+ adc<22> adc<23> adc<24> adc<25> adc<26> adc<27> adc<28> adc<29> adc<30> 
+ adc<31> d<0> d<1> d<2> d<3> d<4> d<5> d<6> d<7> d<8> d<9> d<10> d<11> d<12> 
+ d<13> d<14> d<15> enread q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> 
+ q<10> q<11> q<12> q<13> q<14> q<15> set vdd vss
*.PININFO a_read<0>:I a_read<1>:I a_read<2>:I a_read<3>:I adc<0>:I adc<1>:I 
*.PININFO adc<2>:I adc<3>:I adc<4>:I adc<5>:I adc<6>:I adc<7>:I adc<8>:I 
*.PININFO adc<9>:I adc<10>:I adc<11>:I adc<12>:I adc<13>:I adc<14>:I adc<15>:I 
*.PININFO adc<16>:I adc<17>:I adc<18>:I adc<19>:I adc<20>:I adc<21>:I 
*.PININFO adc<22>:I adc<23>:I adc<24>:I adc<25>:I adc<26>:I adc<27>:I 
*.PININFO adc<28>:I adc<29>:I adc<30>:I adc<31>:I enread:I set:I q<0>:O q<1>:O 
*.PININFO q<2>:O q<3>:O q<4>:O q<5>:O q<6>:O q<7>:O q<8>:O q<9>:O q<10>:O 
*.PININFO q<11>:O q<12>:O q<13>:O q<14>:O q<15>:O d<0>:B d<1>:B d<2>:B d<3>:B 
*.PININFO d<4>:B d<5>:B d<6>:B d<7>:B d<8>:B d<9>:B d<10>:B d<11>:B d<12>:B 
*.PININFO d<13>:B d<14>:B d<15>:B vdd:B vss:B
XI17 adc<30> adc<31> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<15> setn vdd vss / countercell2
XI16 adc<28> adc<29> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<14> setn vdd vss / countercell2
XI15 adc<26> adc<27> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<13> setn vdd vss / countercell2
XI14 adc<24> adc<25> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<12> setn vdd vss / countercell2
XI13 adc<22> adc<23> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<11> setn vdd vss / countercell2
XI12 adc<20> adc<21> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<10> setn vdd vss / countercell2
XI11 adc<18> adc<19> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<9> setn vdd vss / countercell2
XI10 adc<16> adc<17> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<8> setn vdd vss / countercell2
XI9 adc<14> adc<15> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<7> setn vdd vss / countercell2
XI8 adc<12> adc<13> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<6> setn vdd vss / countercell2
XI7 adc<10> adc<11> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> 
+ op<9> op<10> op<11> q<5> setn vdd vss / countercell2
XI6 adc<8> adc<9> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> op<9> 
+ op<10> op<11> q<4> setn vdd vss / countercell2
XI5 adc<6> adc<7> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> op<9> 
+ op<10> op<11> q<3> setn vdd vss / countercell2
XI4 adc<4> adc<5> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> op<9> 
+ op<10> op<11> q<2> setn vdd vss / countercell2
XI3 adc<2> adc<3> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> op<9> 
+ op<10> op<11> q<1> setn vdd vss / countercell2
XI2 adc<0> adc<1> op<0> op<1> op<2> op<3> op<4> op<5> op<6> op<7> op<8> op<9> 
+ op<10> op<11> q<0> setn vdd vss / countercell2
XI20 set setn vdd vss / inv4
XI18 vdd vss enread a_read<0> a_read<1> a_read<2> a_read<3> op<0> op<1> op<2> 
+ op<3> op<4> op<5> net010<0> net010<1> op<6> op<7> op<8> op<9> op<10> op<11> 
+ net011<0> net011<1> / 4x16decoder2
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    invz
* View Name:    schematic
************************************************************************

.SUBCKT invz IN OE OEN OUT VDD VSS
*.PININFO IN:B OE:B OEN:B OUT:B VDD:B VSS:B
XPM3 OUT OEN net13 VDD p12ll_mis_ckt MR=1 L=80n W=200n
XPM2 net13 IN VDD VDD p12ll_mis_ckt MR=1 L=80n W=200n
XNM3 net14 IN VSS VSS n12ll_mis_ckt MR=1 L=80n W=200n
XNM2 OUT OE net14 VSS n12ll_mis_ckt MR=1 L=80n W=200n
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    slatch
* View Name:    schematic
************************************************************************

.SUBCKT slatch clk clkn d q qn vdd vss
*.PININFO clk:I clkn:I d:I q:O qn:O vdd:B vss:B
XI1 net24 clk clkn qn vdd vss / Tgate
XI4 q clkn clk qn vdd vss / invz
XI3 qn q vdd vss / inv2
XI0 d net24 vdd vss / inv2
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    mlatch
* View Name:    schematic
************************************************************************

.SUBCKT mlatch clk clkn d q qn vdd vss
*.PININFO clk:I clkn:I d:I q:O qn:O vdd:B vss:B
XI1 net24 clkn clk qn vdd vss / Tgate
XI4 q clk clkn qn vdd vss / invz
XI3 qn q vdd vss / inv2
XI0 d net24 vdd vss / inv2
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    IO
* View Name:    schematic
************************************************************************

.SUBCKT IO clk_read clk_write d<0> d<1> d<2> d<3> d<4> d<5> d<6> d<7> d<8> 
+ d<9> d<10> d<11> d<12> d<13> d<14> d<15> db<0> db<1> db<2> db<3> db<4> db<5> 
+ db<6> db<7> db<8> db<9> db<10> db<11> db<12> db<13> db<14> db<15> q<0> q<1> 
+ q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> q<14> q<15> 
+ qb<0> qb<1> qb<2> qb<3> qb<4> qb<5> qb<6> qb<7> qb<8> qb<9> qb<10> qb<11> 
+ qb<12> qb<13> qb<14> qb<15> vdd vss
*.PININFO clk_read:I clk_write:I d<0>:I d<1>:I d<2>:I d<3>:I d<4>:I d<5>:I 
*.PININFO d<6>:I d<7>:I d<8>:I d<9>:I d<10>:I d<11>:I d<12>:I d<13>:I d<14>:I 
*.PININFO d<15>:I q<0>:I q<1>:I q<2>:I q<3>:I q<4>:I q<5>:I q<6>:I q<7>:I 
*.PININFO q<8>:I q<9>:I q<10>:I q<11>:I q<12>:I q<13>:I q<14>:I q<15>:I 
*.PININFO db<0>:O db<1>:O db<2>:O db<3>:O db<4>:O db<5>:O db<6>:O db<7>:O 
*.PININFO db<8>:O db<9>:O db<10>:O db<11>:O db<12>:O db<13>:O db<14>:O 
*.PININFO db<15>:O qb<0>:O qb<1>:O qb<2>:O qb<3>:O qb<4>:O qb<5>:O qb<6>:O 
*.PININFO qb<7>:O qb<8>:O qb<9>:O qb<10>:O qb<11>:O qb<12>:O qb<13>:O qb<14>:O 
*.PININFO qb<15>:O vdd:B vss:B
XI8<0> net037<0> net024<0> vdd vss / inv1
XI8<1> net037<1> net024<1> vdd vss / inv1
XI8<2> net037<2> net024<2> vdd vss / inv1
XI8<3> net037<3> net024<3> vdd vss / inv1
XI8<4> net037<4> net024<4> vdd vss / inv1
XI8<5> net037<5> net024<5> vdd vss / inv1
XI8<6> net037<6> net024<6> vdd vss / inv1
XI8<7> net037<7> net024<7> vdd vss / inv1
XI8<8> net037<8> net024<8> vdd vss / inv1
XI8<9> net037<9> net024<9> vdd vss / inv1
XI8<10> net037<10> net024<10> vdd vss / inv1
XI8<11> net037<11> net024<11> vdd vss / inv1
XI8<12> net037<12> net024<12> vdd vss / inv1
XI8<13> net037<13> net024<13> vdd vss / inv1
XI8<14> net037<14> net024<14> vdd vss / inv1
XI8<15> net037<15> net024<15> vdd vss / inv1
XI7<0> q<0> net040<0> vdd vss / inv1
XI7<1> q<1> net040<1> vdd vss / inv1
XI7<2> q<2> net040<2> vdd vss / inv1
XI7<3> q<3> net040<3> vdd vss / inv1
XI7<4> q<4> net040<4> vdd vss / inv1
XI7<5> q<5> net040<5> vdd vss / inv1
XI7<6> q<6> net040<6> vdd vss / inv1
XI7<7> q<7> net040<7> vdd vss / inv1
XI7<8> q<8> net040<8> vdd vss / inv1
XI7<9> q<9> net040<9> vdd vss / inv1
XI7<10> q<10> net040<10> vdd vss / inv1
XI7<11> q<11> net040<11> vdd vss / inv1
XI7<12> q<12> net040<12> vdd vss / inv1
XI7<13> q<13> net040<13> vdd vss / inv1
XI7<14> q<14> net040<14> vdd vss / inv1
XI7<15> q<15> net040<15> vdd vss / inv1
XI6<0> net040<0> net015<0> vdd vss / inv1
XI6<1> net040<1> net015<1> vdd vss / inv1
XI6<2> net040<2> net015<2> vdd vss / inv1
XI6<3> net040<3> net015<3> vdd vss / inv1
XI6<4> net040<4> net015<4> vdd vss / inv1
XI6<5> net040<5> net015<5> vdd vss / inv1
XI6<6> net040<6> net015<6> vdd vss / inv1
XI6<7> net040<7> net015<7> vdd vss / inv1
XI6<8> net040<8> net015<8> vdd vss / inv1
XI6<9> net040<9> net015<9> vdd vss / inv1
XI6<10> net040<10> net015<10> vdd vss / inv1
XI6<11> net040<11> net015<11> vdd vss / inv1
XI6<12> net040<12> net015<12> vdd vss / inv1
XI6<13> net040<13> net015<13> vdd vss / inv1
XI6<14> net040<14> net015<14> vdd vss / inv1
XI6<15> net040<15> net015<15> vdd vss / inv1
XI4<0> net033<0> db<0> vdd vss / inv1
XI4<1> net033<1> db<1> vdd vss / inv1
XI4<2> net033<2> db<2> vdd vss / inv1
XI4<3> net033<3> db<3> vdd vss / inv1
XI4<4> net033<4> db<4> vdd vss / inv1
XI4<5> net033<5> db<5> vdd vss / inv1
XI4<6> net033<6> db<6> vdd vss / inv1
XI4<7> net033<7> db<7> vdd vss / inv1
XI4<8> net033<8> db<8> vdd vss / inv1
XI4<9> net033<9> db<9> vdd vss / inv1
XI4<10> net033<10> db<10> vdd vss / inv1
XI4<11> net033<11> db<11> vdd vss / inv1
XI4<12> net033<12> db<12> vdd vss / inv1
XI4<13> net033<13> db<13> vdd vss / inv1
XI4<14> net033<14> db<14> vdd vss / inv1
XI4<15> net033<15> db<15> vdd vss / inv1
XI3<0> net032<0> net033<0> vdd vss / inv1
XI3<1> net032<1> net033<1> vdd vss / inv1
XI3<2> net032<2> net033<2> vdd vss / inv1
XI3<3> net032<3> net033<3> vdd vss / inv1
XI3<4> net032<4> net033<4> vdd vss / inv1
XI3<5> net032<5> net033<5> vdd vss / inv1
XI3<6> net032<6> net033<6> vdd vss / inv1
XI3<7> net032<7> net033<7> vdd vss / inv1
XI3<8> net032<8> net033<8> vdd vss / inv1
XI3<9> net032<9> net033<9> vdd vss / inv1
XI3<10> net032<10> net033<10> vdd vss / inv1
XI3<11> net032<11> net033<11> vdd vss / inv1
XI3<12> net032<12> net033<12> vdd vss / inv1
XI3<13> net032<13> net033<13> vdd vss / inv1
XI3<14> net032<14> net033<14> vdd vss / inv1
XI3<15> net032<15> net033<15> vdd vss / inv1
XI2<0> net025<0> net016<0> vdd vss / inv1
XI2<1> net025<1> net016<1> vdd vss / inv1
XI2<2> net025<2> net016<2> vdd vss / inv1
XI2<3> net025<3> net016<3> vdd vss / inv1
XI2<4> net025<4> net016<4> vdd vss / inv1
XI2<5> net025<5> net016<5> vdd vss / inv1
XI2<6> net025<6> net016<6> vdd vss / inv1
XI2<7> net025<7> net016<7> vdd vss / inv1
XI2<8> net025<8> net016<8> vdd vss / inv1
XI2<9> net025<9> net016<9> vdd vss / inv1
XI2<10> net025<10> net016<10> vdd vss / inv1
XI2<11> net025<11> net016<11> vdd vss / inv1
XI2<12> net025<12> net016<12> vdd vss / inv1
XI2<13> net025<13> net016<13> vdd vss / inv1
XI2<14> net025<14> net016<14> vdd vss / inv1
XI2<15> net025<15> net016<15> vdd vss / inv1
XI16 clk_read clk_readn vdd vss / inv4
XI15 clk_write clk_writen vdd vss / inv4
XI14 clk_readn clk_readb vdd vss / inv4
XI13 clk_writen clk_writeb vdd vss / inv4
XI12<0> clk_readb clk_readn net017<0> net028<0> net041<0> vdd vss / slatch
XI12<1> clk_readb clk_readn net017<1> net028<1> net041<1> vdd vss / slatch
XI12<2> clk_readb clk_readn net017<2> net028<2> net041<2> vdd vss / slatch
XI12<3> clk_readb clk_readn net017<3> net028<3> net041<3> vdd vss / slatch
XI12<4> clk_readb clk_readn net017<4> net028<4> net041<4> vdd vss / slatch
XI12<5> clk_readb clk_readn net017<5> net028<5> net041<5> vdd vss / slatch
XI12<6> clk_readb clk_readn net017<6> net028<6> net041<6> vdd vss / slatch
XI12<7> clk_readb clk_readn net017<7> net028<7> net041<7> vdd vss / slatch
XI12<8> clk_readb clk_readn net017<8> net028<8> net041<8> vdd vss / slatch
XI12<9> clk_readb clk_readn net017<9> net028<9> net041<9> vdd vss / slatch
XI12<10> clk_readb clk_readn net017<10> net028<10> net041<10> vdd vss / slatch
XI12<11> clk_readb clk_readn net017<11> net028<11> net041<11> vdd vss / slatch
XI12<12> clk_readb clk_readn net017<12> net028<12> net041<12> vdd vss / slatch
XI12<13> clk_readb clk_readn net017<13> net028<13> net041<13> vdd vss / slatch
XI12<14> clk_readb clk_readn net017<14> net028<14> net041<14> vdd vss / slatch
XI12<15> clk_readb clk_readn net017<15> net028<15> net041<15> vdd vss / slatch
XI23<0> clk_writeb clk_writen net029<0> net032<0> net035<0> vdd vss / slatch
XI23<1> clk_writeb clk_writen net029<1> net032<1> net035<1> vdd vss / slatch
XI23<2> clk_writeb clk_writen net029<2> net032<2> net035<2> vdd vss / slatch
XI23<3> clk_writeb clk_writen net029<3> net032<3> net035<3> vdd vss / slatch
XI23<4> clk_writeb clk_writen net029<4> net032<4> net035<4> vdd vss / slatch
XI23<5> clk_writeb clk_writen net029<5> net032<5> net035<5> vdd vss / slatch
XI23<6> clk_writeb clk_writen net029<6> net032<6> net035<6> vdd vss / slatch
XI23<7> clk_writeb clk_writen net029<7> net032<7> net035<7> vdd vss / slatch
XI23<8> clk_writeb clk_writen net029<8> net032<8> net035<8> vdd vss / slatch
XI23<9> clk_writeb clk_writen net029<9> net032<9> net035<9> vdd vss / slatch
XI23<10> clk_writeb clk_writen net029<10> net032<10> net035<10> vdd vss / 
+ slatch
XI23<11> clk_writeb clk_writen net029<11> net032<11> net035<11> vdd vss / 
+ slatch
XI23<12> clk_writeb clk_writen net029<12> net032<12> net035<12> vdd vss / 
+ slatch
XI23<13> clk_writeb clk_writen net029<13> net032<13> net035<13> vdd vss / 
+ slatch
XI23<14> clk_writeb clk_writen net029<14> net032<14> net035<14> vdd vss / 
+ slatch
XI23<15> clk_writeb clk_writen net029<15> net032<15> net035<15> vdd vss / 
+ slatch
XI11<0> clk_readb clk_readn net028<0> net037<0> net039<0> vdd vss / mlatch
XI11<1> clk_readb clk_readn net028<1> net037<1> net039<1> vdd vss / mlatch
XI11<2> clk_readb clk_readn net028<2> net037<2> net039<2> vdd vss / mlatch
XI11<3> clk_readb clk_readn net028<3> net037<3> net039<3> vdd vss / mlatch
XI11<4> clk_readb clk_readn net028<4> net037<4> net039<4> vdd vss / mlatch
XI11<5> clk_readb clk_readn net028<5> net037<5> net039<5> vdd vss / mlatch
XI11<6> clk_readb clk_readn net028<6> net037<6> net039<6> vdd vss / mlatch
XI11<7> clk_readb clk_readn net028<7> net037<7> net039<7> vdd vss / mlatch
XI11<8> clk_readb clk_readn net028<8> net037<8> net039<8> vdd vss / mlatch
XI11<9> clk_readb clk_readn net028<9> net037<9> net039<9> vdd vss / mlatch
XI11<10> clk_readb clk_readn net028<10> net037<10> net039<10> vdd vss / mlatch
XI11<11> clk_readb clk_readn net028<11> net037<11> net039<11> vdd vss / mlatch
XI11<12> clk_readb clk_readn net028<12> net037<12> net039<12> vdd vss / mlatch
XI11<13> clk_readb clk_readn net028<13> net037<13> net039<13> vdd vss / mlatch
XI11<14> clk_readb clk_readn net028<14> net037<14> net039<14> vdd vss / mlatch
XI11<15> clk_readb clk_readn net028<15> net037<15> net039<15> vdd vss / mlatch
XI24<0> clk_writeb clk_writen net018<0> net029<0> net036<0> vdd vss / mlatch
XI24<1> clk_writeb clk_writen net018<1> net029<1> net036<1> vdd vss / mlatch
XI24<2> clk_writeb clk_writen net018<2> net029<2> net036<2> vdd vss / mlatch
XI24<3> clk_writeb clk_writen net018<3> net029<3> net036<3> vdd vss / mlatch
XI24<4> clk_writeb clk_writen net018<4> net029<4> net036<4> vdd vss / mlatch
XI24<5> clk_writeb clk_writen net018<5> net029<5> net036<5> vdd vss / mlatch
XI24<6> clk_writeb clk_writen net018<6> net029<6> net036<6> vdd vss / mlatch
XI24<7> clk_writeb clk_writen net018<7> net029<7> net036<7> vdd vss / mlatch
XI24<8> clk_writeb clk_writen net018<8> net029<8> net036<8> vdd vss / mlatch
XI24<9> clk_writeb clk_writen net018<9> net029<9> net036<9> vdd vss / mlatch
XI24<10> clk_writeb clk_writen net018<10> net029<10> net036<10> vdd vss / 
+ mlatch
XI24<11> clk_writeb clk_writen net018<11> net029<11> net036<11> vdd vss / 
+ mlatch
XI24<12> clk_writeb clk_writen net018<12> net029<12> net036<12> vdd vss / 
+ mlatch
XI24<13> clk_writeb clk_writen net018<13> net029<13> net036<13> vdd vss / 
+ mlatch
XI24<14> clk_writeb clk_writen net018<14> net029<14> net036<14> vdd vss / 
+ mlatch
XI24<15> clk_writeb clk_writen net018<15> net029<15> net036<15> vdd vss / 
+ mlatch
XI9<0> net024<0> qb<0> vdd vss / inv8
XI9<1> net024<1> qb<1> vdd vss / inv8
XI9<2> net024<2> qb<2> vdd vss / inv8
XI9<3> net024<3> qb<3> vdd vss / inv8
XI9<4> net024<4> qb<4> vdd vss / inv8
XI9<5> net024<5> qb<5> vdd vss / inv8
XI9<6> net024<6> qb<6> vdd vss / inv8
XI9<7> net024<7> qb<7> vdd vss / inv8
XI9<8> net024<8> qb<8> vdd vss / inv8
XI9<9> net024<9> qb<9> vdd vss / inv8
XI9<10> net024<10> qb<10> vdd vss / inv8
XI9<11> net024<11> qb<11> vdd vss / inv8
XI9<12> net024<12> qb<12> vdd vss / inv8
XI9<13> net024<13> qb<13> vdd vss / inv8
XI9<14> net024<14> qb<14> vdd vss / inv8
XI9<15> net024<15> qb<15> vdd vss / inv8
XI20<0> d<0> net025<0> vdd vss / inv8
XI20<1> d<1> net025<1> vdd vss / inv8
XI20<2> d<2> net025<2> vdd vss / inv8
XI20<3> d<3> net025<3> vdd vss / inv8
XI20<4> d<4> net025<4> vdd vss / inv8
XI20<5> d<5> net025<5> vdd vss / inv8
XI20<6> d<6> net025<6> vdd vss / inv8
XI20<7> d<7> net025<7> vdd vss / inv8
XI20<8> d<8> net025<8> vdd vss / inv8
XI20<9> d<9> net025<9> vdd vss / inv8
XI20<10> d<10> net025<10> vdd vss / inv8
XI20<11> d<11> net025<11> vdd vss / inv8
XI20<12> d<12> net025<12> vdd vss / inv8
XI20<13> d<13> net025<13> vdd vss / inv8
XI20<14> d<14> net025<14> vdd vss / inv8
XI20<15> d<15> net025<15> vdd vss / inv8
XI19<0> vdd vss net016<0> net018<0> / delaycell_editable
XI19<1> vdd vss net016<1> net018<1> / delaycell_editable
XI19<2> vdd vss net016<2> net018<2> / delaycell_editable
XI19<3> vdd vss net016<3> net018<3> / delaycell_editable
XI19<4> vdd vss net016<4> net018<4> / delaycell_editable
XI19<5> vdd vss net016<5> net018<5> / delaycell_editable
XI19<6> vdd vss net016<6> net018<6> / delaycell_editable
XI19<7> vdd vss net016<7> net018<7> / delaycell_editable
XI19<8> vdd vss net016<8> net018<8> / delaycell_editable
XI19<9> vdd vss net016<9> net018<9> / delaycell_editable
XI19<10> vdd vss net016<10> net018<10> / delaycell_editable
XI19<11> vdd vss net016<11> net018<11> / delaycell_editable
XI19<12> vdd vss net016<12> net018<12> / delaycell_editable
XI19<13> vdd vss net016<13> net018<13> / delaycell_editable
XI19<14> vdd vss net016<14> net018<14> / delaycell_editable
XI19<15> vdd vss net016<15> net018<15> / delaycell_editable
XI21<0> vdd vss net015<0> net017<0> / delaycell_editable
XI21<1> vdd vss net015<1> net017<1> / delaycell_editable
XI21<2> vdd vss net015<2> net017<2> / delaycell_editable
XI21<3> vdd vss net015<3> net017<3> / delaycell_editable
XI21<4> vdd vss net015<4> net017<4> / delaycell_editable
XI21<5> vdd vss net015<5> net017<5> / delaycell_editable
XI21<6> vdd vss net015<6> net017<6> / delaycell_editable
XI21<7> vdd vss net015<7> net017<7> / delaycell_editable
XI21<8> vdd vss net015<8> net017<8> / delaycell_editable
XI21<9> vdd vss net015<9> net017<9> / delaycell_editable
XI21<10> vdd vss net015<10> net017<10> / delaycell_editable
XI21<11> vdd vss net015<11> net017<11> / delaycell_editable
XI21<12> vdd vss net015<12> net017<12> / delaycell_editable
XI21<13> vdd vss net015<13> net017<13> / delaycell_editable
XI21<14> vdd vss net015<14> net017<14> / delaycell_editable
XI21<15> vdd vss net015<15> net017<15> / delaycell_editable
.ENDS

************************************************************************
* Library Name: LogicGates
* Cell Name:    Tgate2
* View Name:    schematic
************************************************************************

.SUBCKT Tgate2 IN OE OEN OUT VDD VSS
*.PININFO IN:B OE:B OEN:B OUT:B VDD:B VSS:B
XNM2 OUT OE IN VSS n12ll_mis_ckt MR=1 L=80n W=600n
XPM0 IN OEN OUT VDD p12ll_mis_ckt MR=1 L=80n W=600n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    SA2
* View Name:    schematic
************************************************************************

.SUBCKT SA2 in1 in2 out vb vdd vss
*.PININFO in1:I in2:I vb:I vdd:I vss:I out:B
XNM8 net015 net015 vss vss n12ll_mis_ckt MR=1 L=80n W=150n
XNM0 net01 net015 vss vss n12ll_mis_ckt MR=1 L=80n W=150n
XNM7 net07 net015 vss vss n12ll_mis_ckt MR=1 L=80n W=300n
XNM9 out net01 vss vss n12ll_mis_ckt MR=1 L=80n W=300n
XPM7 net07 net07 vdd vdd p12ll_mis_ckt MR=1 L=80n W=600n
XPM5 net01 in2 net26 vdd p12ll_mis_ckt MR=1 L=80n W=300n
XPM4 net26 vb vdd vdd p12ll_mis_ckt MR=1 L=80n W=300n
XPM8 net015 in1 net26 vdd p12ll_mis_ckt MR=1 L=80n W=300n
XPM9 out net07 vdd vdd p12ll_mis_ckt MR=1 L=80n W=600n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    ADCcell
* View Name:    schematic
************************************************************************

.SUBCKT ADCcell cbl model modeln set set_comp set_compn setn vb vb2 vb3 vdd 
+ vss x<5>
*.PININFO cbl:I model:I modeln:I set:I set_comp:I set_compn:I setn:I vb:I 
*.PININFO vb2:I vb3:I vdd:I vss:I x<5>:O
XI23 net54 net014 vdd vss / inv0_5
XI22 x<1> set net54 vdd vss / nor
XNM5 Vc x<3> vss vss n12ll_mis_ckt MR=1 L=80n W=1.2u
XNM4 vss set_compn x<1> vss n12ll_mis_ckt MR=1 L=80n W=300n
XNM3 net016 bc Vc vss n12ll_mis_ckt MR=1 L=80n W=1.2u
XNM2 cbl vb3 net016 vss n12ll_mis_ckt MR=1 L=80n W=600n
XNM6 Vc set vss vss n12ll_mis_ckt MR=1 L=80n W=600n
XI7 x<0> set_comp set_compn x<1> vdd vss / invz
XI1 cbl set setn vb vdd vss / Tgate
XI3<0> x<1> x<2> vdd vss / inv0_3
XI3<1> x<2> x<3> vdd vss / inv0_3
XI3<2> x<3> x<4> vdd vss / inv0_3
XI4 Vc modeln model net010 vdd vss / Tgate2
XI8 x<4> x<5> vdd vss / inv1
XI5 net014 bc vdd vss / inv1
XI0 Vc vb x<0> vb2 vdd vss / SA2
XC0 net010 vss mom_2t_ckt LF=5.3u NF=22 TM=3 BM=1 MR=1
XC2 cbl vss mom_2t_ckt LF=10u NF=20 TM=3 BM=1 MR=1
XC1 Vc vss mom_2t_ckt LF=5.3u NF=5 TM=3 BM=1 MR=1
XPM0 vdd set_comp vb2 vdd p12ll_mis_ckt MR=1 L=80n W=1.2u
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    SA
* View Name:    schematic
************************************************************************

.SUBCKT SA in1 in2 out vb vdd vss
*.PININFO in1:I in2:I vb:I out:B vdd:B vss:B
XPM2 net021 in2 net16 vdd p12ll_mis_ckt MR=1 L=120n W=600n
XPM3 net019 in1 net16 vdd p12ll_mis_ckt MR=1 L=120n W=600n
XPM0 net07 net07 vdd vdd p12ll_mis_ckt MR=1 L=120n W=2.4u
XPM1 net16 vb vdd vdd p12ll_mis_ckt MR=1 L=120n W=600n
XPM4 out net07 vdd vdd p12ll_mis_ckt MR=1 L=120n W=19.2u
XNM1 net07 net019 vss vss n12ll_mis_ckt MR=1 L=120n W=1.2u
XNM2 net021 net019 vss vss n12ll_mis_ckt MR=1 L=120n W=300n
XNM3 out net021 vss vss n12ll_mis_ckt MR=1 L=120n W=9.6u
XNM0 net019 net019 vss vss n12ll_mis_ckt MR=1 L=120n W=300n
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    bias
* View Name:    schematic
************************************************************************

.SUBCKT bias set set_comp vb vb2 vb3 vdd vss
*.PININFO set:I set_comp:I vb:O vb2:O vb3:O vdd:B vss:B
RR7 vdd net028 70.5375K $[rnwsti] $W=1.6u $L=150u M=1
RR6 vdd net011 70.5375K $[rnwsti] $W=1.6u $L=150u M=1
RR8 vdd net027 94.05K $[rnwsti] $W=1.6u $L=200u M=1
RR9 vdd net05 94.05K $[rnwsti] $W=1.6u $L=200u M=1
XI36 net010 setn setb vb vdd vss / Tgate
XI38 vb2 setb setn net09 vdd vss / Tgate
XI37 net018 setb setn vb vdd vss / Tgate
XI39 vbr set_compb set_compn net010 vdd vss / Tgate
XI35 setn setb vdd vss / inv4
XI34 set setn vdd vss / inv4
XI10 set_compn set_compb vdd vss / inv4
XI9 set_comp set_compn vdd vss / inv4
XI25 vb net010 net018 net09 vdd vss / SA
XPM0 vbr vbr vdd vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM2 vb3 set_compn net05 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM6 vb3 set_compn net027 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM7 vb2 set_compn net011 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM9 vb2 set_compn net028 vdd p12ll_mis_ckt MR=1 L=600n W=1u
XPM10 net09 setb vdd vdd p12ll_mis_ckt MR=1 L=600n W=600n
XPM1 vbr vbr vdd vdd p12ll_mis_ckt MR=1 L=600n W=1u
XNM6 vbr set_compb net026 vss n12ll_mis_ckt MR=1 L=600n W=1u
XNM15 vb2 vb2 vss vss n12ll_mis_ckt MR=1 L=600n W=500n
XNM16 vbr set_compb net1 vss n12ll_mis_ckt MR=1 L=600n W=1u
XNM10 vb3 vb3 vss vss n12ll_mis_ckt MR=1 L=600n W=600n
XNM12 vb2 vb2 vss vss n12ll_mis_ckt MR=1 L=600n W=500n
XNM11 vb3 vb3 vss vss n12ll_mis_ckt MR=1 L=600n W=600n
XR0 net026 vss rhrpo_ckt M=1 W=7u L=30u
XR1 net1 vss rhrpo_ckt M=1 W=7u L=30u
XC8 vb2 vss mom_2t_ckt LF=30u NF=52 TM=3 BM=1 MR=1
XC9 vb vss mom_2t_ckt LF=30u NF=52 TM=3 BM=1 MR=1
XC5 vb3 vss mom_2t_ckt LF=30u NF=52 TM=3 BM=1 MR=1
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    ADC
* View Name:    schematic
************************************************************************

.SUBCKT ADC adc<0> adc<1> adc<2> adc<3> adc<4> adc<5> adc<6> adc<7> adc<8> 
+ adc<9> adc<10> adc<11> adc<12> adc<13> adc<14> adc<15> adc<16> adc<17> 
+ adc<18> adc<19> adc<20> adc<21> adc<22> adc<23> adc<24> adc<25> adc<26> 
+ adc<27> adc<28> adc<29> adc<30> adc<31> cbl<0> cbl<1> cbl<2> cbl<3> cbl<4> 
+ cbl<5> cbl<6> cbl<7> cbl<8> cbl<9> cbl<10> cbl<11> cbl<12> cbl<13> cbl<14> 
+ cbl<15> cbl<16> cbl<17> cbl<18> cbl<19> cbl<20> cbl<21> cbl<22> cbl<23> 
+ cbl<24> cbl<25> cbl<26> cbl<27> cbl<28> cbl<29> cbl<30> cbl<31> d<0> d<1> 
+ d<2> d<3> d<4> d<5> d<6> d<7> d<8> d<9> d<10> d<11> d<12> d<13> d<14> d<15> 
+ model set set_comp vdd vss
*.PININFO cbl<0>:I cbl<1>:I cbl<2>:I cbl<3>:I cbl<4>:I cbl<5>:I cbl<6>:I 
*.PININFO cbl<7>:I cbl<8>:I cbl<9>:I cbl<10>:I cbl<11>:I cbl<12>:I cbl<13>:I 
*.PININFO cbl<14>:I cbl<15>:I cbl<16>:I cbl<17>:I cbl<18>:I cbl<19>:I 
*.PININFO cbl<20>:I cbl<21>:I cbl<22>:I cbl<23>:I cbl<24>:I cbl<25>:I 
*.PININFO cbl<26>:I cbl<27>:I cbl<28>:I cbl<29>:I cbl<30>:I cbl<31>:I model:I 
*.PININFO set:I set_comp:I adc<0>:O adc<1>:O adc<2>:O adc<3>:O adc<4>:O 
*.PININFO adc<5>:O adc<6>:O adc<7>:O adc<8>:O adc<9>:O adc<10>:O adc<11>:O 
*.PININFO adc<12>:O adc<13>:O adc<14>:O adc<15>:O adc<16>:O adc<17>:O 
*.PININFO adc<18>:O adc<19>:O adc<20>:O adc<21>:O adc<22>:O adc<23>:O 
*.PININFO adc<24>:O adc<25>:O adc<26>:O adc<27>:O adc<28>:O adc<29>:O 
*.PININFO adc<30>:O adc<31>:O d<0>:B d<1>:B d<2>:B d<3>:B d<4>:B d<5>:B d<6>:B 
*.PININFO d<7>:B d<8>:B d<9>:B d<10>:B d<11>:B d<12>:B d<13>:B d<14>:B d<15>:B 
*.PININFO vdd:B vss:B
XI0<0> cbl<0> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<0> / ADCcell
XI0<1> cbl<1> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<1> / ADCcell
XI0<2> cbl<2> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<2> / ADCcell
XI0<3> cbl<3> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<3> / ADCcell
XI0<4> cbl<4> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<4> / ADCcell
XI0<5> cbl<5> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<5> / ADCcell
XI0<6> cbl<6> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<6> / ADCcell
XI0<7> cbl<7> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<7> / ADCcell
XI0<8> cbl<8> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<8> / ADCcell
XI0<9> cbl<9> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd vss 
+ adc<9> / ADCcell
XI0<10> cbl<10> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<10> / ADCcell
XI0<11> cbl<11> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<11> / ADCcell
XI0<12> cbl<12> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<12> / ADCcell
XI0<13> cbl<13> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<13> / ADCcell
XI0<14> cbl<14> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<14> / ADCcell
XI0<15> cbl<15> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<15> / ADCcell
XI0<16> cbl<16> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<16> / ADCcell
XI0<17> cbl<17> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<17> / ADCcell
XI0<18> cbl<18> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<18> / ADCcell
XI0<19> cbl<19> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<19> / ADCcell
XI0<20> cbl<20> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<20> / ADCcell
XI0<21> cbl<21> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<21> / ADCcell
XI0<22> cbl<22> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<22> / ADCcell
XI0<23> cbl<23> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<23> / ADCcell
XI0<24> cbl<24> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<24> / ADCcell
XI0<25> cbl<25> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<25> / ADCcell
XI0<26> cbl<26> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<26> / ADCcell
XI0<27> cbl<27> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<27> / ADCcell
XI0<28> cbl<28> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<28> / ADCcell
XI0<29> cbl<29> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<29> / ADCcell
XI0<30> cbl<30> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<30> / ADCcell
XI0<31> cbl<31> modelb modelbn setb set_compb set_compn setbn vb vb2 vb3 vdd 
+ vss adc<31> / ADCcell
XI7 set_compn set_compb vdd vss / inv4
XI6 set_comp set_compn vdd vss / inv4
XI3 modelbn modelb vdd vss / inv4
XI2 model modelbn vdd vss / inv4
XI1 setbn setb vdd vss / inv4
XI16 set setbn vdd vss / inv4
XI5 setb set_compb vb vb2 vb3 vdd vss / bias
.ENDS

************************************************************************
* Library Name: SRAM_ChargePulsation
* Cell Name:    SRAM_CIM
* View Name:    schematic
************************************************************************

.SUBCKT SRAM_CIM a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> clk comp d<15> 
+ d<14> d<13> d<12> d<11> d<10> d<9> d<8> d<7> d<6> d<5> d<4> d<3> d<2> d<1> 
+ d<0> inbit model q<15> q<14> q<13> q<12> q<11> q<10> q<9> q<8> q<7> q<6> q<5> 
+ q<4> q<3> q<2> q<1> q<0> read set wait_ wrt wrtbuf
*.PININFO a<0>:I a<1>:I a<2>:I a<3>:I a<4>:I a<5>:I a<6>:I a<7>:I a<8>:I clk:I 
*.PININFO comp:I d<0>:I d<1>:I d<2>:I d<3>:I d<4>:I d<5>:I d<6>:I d<7>:I 
*.PININFO d<8>:I d<9>:I d<10>:I d<11>:I d<12>:I d<13>:I d<14>:I d<15>:I 
*.PININFO inbit:I model:I read:I set:I wait_:I wrt:I wrtbuf:I q<0>:O q<1>:O 
*.PININFO q<2>:O q<3>:O q<4>:O q<5>:O q<6>:O q<7>:O q<8>:O q<9>:O q<10>:O 
*.PININFO q<11>:O q<12>:O q<13>:O q<14>:O q<15>:O vdd:B vss:B
XI0 net8<0> net8<1> net8<2> net8<3> net8<4> net8<5> net8<6> net8<7> net8<8> 
+ net8<9> net8<10> net8<11> net8<12> net8<13> net8<14> net8<15> net8<16> 
+ net8<17> net8<18> net8<19> net8<20> net8<21> net8<22> net8<23> net8<24> 
+ net8<25> net8<26> net8<27> net8<28> net8<29> net8<30> net8<31> net8<32> 
+ net8<33> net8<34> net8<35> net8<36> net8<37> net8<38> net8<39> net8<40> 
+ net8<41> net8<42> net8<43> net8<44> net8<45> net8<46> net8<47> net8<48> 
+ net8<49> net8<50> net8<51> net8<52> net8<53> net8<54> net8<55> net8<56> 
+ net8<57> net8<58> net8<59> net8<60> net8<61> net8<62> net8<63> net035<0> 
+ net035<1> net035<2> net035<3> net035<4> net035<5> net035<6> net035<7> 
+ net035<8> net035<9> net035<10> net035<11> net035<12> net035<13> net035<14> 
+ net035<15> net072<0> net072<1> net072<2> net072<3> net072<4> net072<5> 
+ net072<6> net072<7> net072<8> net072<9> net072<10> net072<11> net072<12> 
+ net072<13> net072<14> net072<15> net072<16> net072<17> net072<18> net072<19> 
+ net072<20> net072<21> net072<22> net072<23> net072<24> net072<25> net072<26> 
+ net072<27> net072<28> net072<29> net072<30> net072<31> net4<0> net4<1> 
+ net4<2> net4<3> net4<4> net4<5> net4<6> net4<7> net4<8> net4<9> net4<10> 
+ net4<11> net4<12> net4<13> net4<14> net4<15> net4<16> net4<17> net4<18> 
+ net4<19> net4<20> net4<21> net4<22> net4<23> net4<24> net4<25> net4<26> 
+ net4<27> net4<28> net4<29> net4<30> net4<31> net4<32> net4<33> net4<34> 
+ net4<35> net4<36> net4<37> net4<38> net4<39> net4<40> net4<41> net4<42> 
+ net4<43> net4<44> net4<45> net4<46> net4<47> net4<48> net4<49> net4<50> 
+ net4<51> net4<52> net4<53> net4<54> net4<55> net4<56> net4<57> net4<58> 
+ net4<59> net4<60> net4<61> net4<62> net4<63> net4<64> net4<65> net4<66> 
+ net4<67> net4<68> net4<69> net4<70> net4<71> net4<72> net4<73> net4<74> 
+ net4<75> net4<76> net4<77> net4<78> net4<79> net4<80> net4<81> net4<82> 
+ net4<83> net4<84> net4<85> net4<86> net4<87> net4<88> net4<89> net4<90> 
+ net4<91> net4<92> net4<93> net4<94> net4<95> net4<96> net4<97> net4<98> 
+ net4<99> net4<100> net4<101> net4<102> net4<103> net4<104> net4<105> 
+ net4<106> net4<107> net4<108> net4<109> net4<110> net4<111> net4<112> 
+ net4<113> net4<114> net4<115> net4<116> net4<117> net4<118> net4<119> 
+ net4<120> net4<121> net4<122> net4<123> net4<124> net4<125> net4<126> 
+ net4<127> net5<0> net5<1> net5<2> net5<3> net5<4> net5<5> net5<6> net5<7> 
+ net5<8> net5<9> net5<10> net5<11> net5<12> net5<13> net5<14> net5<15> 
+ net5<16> net5<17> net5<18> net5<19> net5<20> net5<21> net5<22> net5<23> 
+ net5<24> net5<25> net5<26> net5<27> net5<28> net5<29> net5<30> net5<31> 
+ net5<32> net5<33> net5<34> net5<35> net5<36> net5<37> net5<38> net5<39> 
+ net5<40> net5<41> net5<42> net5<43> net5<44> net5<45> net5<46> net5<47> 
+ net5<48> net5<49> net5<50> net5<51> net5<52> net5<53> net5<54> net5<55> 
+ net5<56> net5<57> net5<58> net5<59> net5<60> net5<61> net5<62> net5<63> 
+ net5<64> net5<65> net5<66> net5<67> net5<68> net5<69> net5<70> net5<71> 
+ net5<72> net5<73> net5<74> net5<75> net5<76> net5<77> net5<78> net5<79> 
+ net5<80> net5<81> net5<82> net5<83> net5<84> net5<85> net5<86> net5<87> 
+ net5<88> net5<89> net5<90> net5<91> net5<92> net5<93> net5<94> net5<95> 
+ net5<96> net5<97> net5<98> net5<99> net5<100> net5<101> net5<102> net5<103> 
+ net5<104> net5<105> net5<106> net5<107> net5<108> net5<109> net5<110> 
+ net5<111> net5<112> net5<113> net5<114> net5<115> net5<116> net5<117> 
+ net5<118> net5<119> net5<120> net5<121> net5<122> net5<123> net5<124> 
+ net5<125> net5<126> net5<127> net6<0> net6<1> net6<2> net6<3> net6<4> 
+ net6<5> net6<6> net6<7> net6<8> net6<9> net6<10> net6<11> net6<12> net6<13> 
+ net6<14> net6<15> net6<16> net6<17> net6<18> net6<19> net6<20> net6<21> 
+ net6<22> net6<23> net6<24> net6<25> net6<26> net6<27> net6<28> net6<29> 
+ net6<30> net6<31> net6<32> net6<33> net6<34> net6<35> net6<36> net6<37> 
+ net6<38> net6<39> net6<40> net6<41> net6<42> net6<43> net6<44> net6<45> 
+ net6<46> net6<47> net6<48> net6<49> net6<50> net6<51> net6<52> net6<53> 
+ net6<54> net6<55> net6<56> net6<57> net6<58> net6<59> net6<60> net6<61> 
+ net6<62> net6<63> net036<0> net036<1> net036<2> net036<3> net036<4> 
+ net036<5> net036<6> net036<7> net036<8> net036<9> net036<10> net036<11> 
+ net036<12> net036<13> net036<14> net036<15> vdd vss net1<0> net1<1> net1<2> 
+ net1<3> net1<4> net1<5> net1<6> net1<7> net1<8> net1<9> net1<10> net1<11> 
+ net1<12> net1<13> net1<14> net1<15> net1<16> net1<17> net1<18> net1<19> 
+ net1<20> net1<21> net1<22> net1<23> net1<24> net1<25> net1<26> net1<27> 
+ net1<28> net1<29> net1<30> net1<31> net1<32> net1<33> net1<34> net1<35> 
+ net1<36> net1<37> net1<38> net1<39> net1<40> net1<41> net1<42> net1<43> 
+ net1<44> net1<45> net1<46> net1<47> net1<48> net1<49> net1<50> net1<51> 
+ net1<52> net1<53> net1<54> net1<55> net1<56> net1<57> net1<58> net1<59> 
+ net1<60> net1<61> net1<62> net1<63> net1<64> net1<65> net1<66> net1<67> 
+ net1<68> net1<69> net1<70> net1<71> net1<72> net1<73> net1<74> net1<75> 
+ net1<76> net1<77> net1<78> net1<79> net1<80> net1<81> net1<82> net1<83> 
+ net1<84> net1<85> net1<86> net1<87> net1<88> net1<89> net1<90> net1<91> 
+ net1<92> net1<93> net1<94> net1<95> net1<96> net1<97> net1<98> net1<99> 
+ net1<100> net1<101> net1<102> net1<103> net1<104> net1<105> net1<106> 
+ net1<107> net1<108> net1<109> net1<110> net1<111> net1<112> net1<113> 
+ net1<114> net1<115> net1<116> net1<117> net1<118> net1<119> net1<120> 
+ net1<121> net1<122> net1<123> net1<124> net1<125> net1<126> net1<127> / array
XI1 net035<0> net035<1> net035<2> net035<3> net035<4> net035<5> net035<6> 
+ net035<7> net035<8> net035<9> net035<10> net035<11> net035<12> net035<13> 
+ net035<14> net035<15> net10<0> net10<1> net10<2> net10<3> net10<4> net10<5> 
+ net10<6> net10<7> net4<0> net4<1> net4<2> net4<3> net4<4> net4<5> net4<6> 
+ net4<7> net4<8> net4<9> net4<10> net4<11> net4<12> net4<13> net4<14> 
+ net4<15> net4<16> net4<17> net4<18> net4<19> net4<20> net4<21> net4<22> 
+ net4<23> net4<24> net4<25> net4<26> net4<27> net4<28> net4<29> net4<30> 
+ net4<31> net4<32> net4<33> net4<34> net4<35> net4<36> net4<37> net4<38> 
+ net4<39> net4<40> net4<41> net4<42> net4<43> net4<44> net4<45> net4<46> 
+ net4<47> net4<48> net4<49> net4<50> net4<51> net4<52> net4<53> net4<54> 
+ net4<55> net4<56> net4<57> net4<58> net4<59> net4<60> net4<61> net4<62> 
+ net4<63> net4<64> net4<65> net4<66> net4<67> net4<68> net4<69> net4<70> 
+ net4<71> net4<72> net4<73> net4<74> net4<75> net4<76> net4<77> net4<78> 
+ net4<79> net4<80> net4<81> net4<82> net4<83> net4<84> net4<85> net4<86> 
+ net4<87> net4<88> net4<89> net4<90> net4<91> net4<92> net4<93> net4<94> 
+ net4<95> net4<96> net4<97> net4<98> net4<99> net4<100> net4<101> net4<102> 
+ net4<103> net4<104> net4<105> net4<106> net4<107> net4<108> net4<109> 
+ net4<110> net4<111> net4<112> net4<113> net4<114> net4<115> net4<116> 
+ net4<117> net4<118> net4<119> net4<120> net4<121> net4<122> net4<123> 
+ net4<124> net4<125> net4<126> net4<127> net5<0> net5<1> net5<2> net5<3> 
+ net5<4> net5<5> net5<6> net5<7> net5<8> net5<9> net5<10> net5<11> net5<12> 
+ net5<13> net5<14> net5<15> net5<16> net5<17> net5<18> net5<19> net5<20> 
+ net5<21> net5<22> net5<23> net5<24> net5<25> net5<26> net5<27> net5<28> 
+ net5<29> net5<30> net5<31> net5<32> net5<33> net5<34> net5<35> net5<36> 
+ net5<37> net5<38> net5<39> net5<40> net5<41> net5<42> net5<43> net5<44> 
+ net5<45> net5<46> net5<47> net5<48> net5<49> net5<50> net5<51> net5<52> 
+ net5<53> net5<54> net5<55> net5<56> net5<57> net5<58> net5<59> net5<60> 
+ net5<61> net5<62> net5<63> net5<64> net5<65> net5<66> net5<67> net5<68> 
+ net5<69> net5<70> net5<71> net5<72> net5<73> net5<74> net5<75> net5<76> 
+ net5<77> net5<78> net5<79> net5<80> net5<81> net5<82> net5<83> net5<84> 
+ net5<85> net5<86> net5<87> net5<88> net5<89> net5<90> net5<91> net5<92> 
+ net5<93> net5<94> net5<95> net5<96> net5<97> net5<98> net5<99> net5<100> 
+ net5<101> net5<102> net5<103> net5<104> net5<105> net5<106> net5<107> 
+ net5<108> net5<109> net5<110> net5<111> net5<112> net5<113> net5<114> 
+ net5<115> net5<116> net5<117> net5<118> net5<119> net5<120> net5<121> 
+ net5<122> net5<123> net5<124> net5<125> net5<126> net5<127> net9<0> net9<1> 
+ net9<2> net9<3> net9<4> net9<5> net9<6> net9<7> net9<8> net9<9> net9<10> 
+ net9<11> net9<12> net9<13> net9<14> net9<15> net036<0> net036<1> net036<2> 
+ net036<3> net036<4> net036<5> net036<6> net036<7> net036<8> net036<9> 
+ net036<10> net036<11> net036<12> net036<13> net036<14> net036<15> vdd vss 
+ net1<0> net1<1> net1<2> net1<3> net1<4> net1<5> net1<6> net1<7> net1<8> 
+ net1<9> net1<10> net1<11> net1<12> net1<13> net1<14> net1<15> net1<16> 
+ net1<17> net1<18> net1<19> net1<20> net1<21> net1<22> net1<23> net1<24> 
+ net1<25> net1<26> net1<27> net1<28> net1<29> net1<30> net1<31> net1<32> 
+ net1<33> net1<34> net1<35> net1<36> net1<37> net1<38> net1<39> net1<40> 
+ net1<41> net1<42> net1<43> net1<44> net1<45> net1<46> net1<47> net1<48> 
+ net1<49> net1<50> net1<51> net1<52> net1<53> net1<54> net1<55> net1<56> 
+ net1<57> net1<58> net1<59> net1<60> net1<61> net1<62> net1<63> net1<64> 
+ net1<65> net1<66> net1<67> net1<68> net1<69> net1<70> net1<71> net1<72> 
+ net1<73> net1<74> net1<75> net1<76> net1<77> net1<78> net1<79> net1<80> 
+ net1<81> net1<82> net1<83> net1<84> net1<85> net1<86> net1<87> net1<88> 
+ net1<89> net1<90> net1<91> net1<92> net1<93> net1<94> net1<95> net1<96> 
+ net1<97> net1<98> net1<99> net1<100> net1<101> net1<102> net1<103> net1<104> 
+ net1<105> net1<106> net1<107> net1<108> net1<109> net1<110> net1<111> 
+ net1<112> net1<113> net1<114> net1<115> net1<116> net1<117> net1<118> 
+ net1<119> net1<120> net1<121> net1<122> net1<123> net1<124> net1<125> 
+ net1<126> net1<127> / WLdriver
XI2 net8<0> net8<1> net8<2> net8<3> net8<4> net8<5> net8<6> net8<7> net8<8> 
+ net8<9> net8<10> net8<11> net8<12> net8<13> net8<14> net8<15> net8<16> 
+ net8<17> net8<18> net8<19> net8<20> net8<21> net8<22> net8<23> net8<24> 
+ net8<25> net8<26> net8<27> net8<28> net8<29> net8<30> net8<31> net8<32> 
+ net8<33> net8<34> net8<35> net8<36> net8<37> net8<38> net8<39> net8<40> 
+ net8<41> net8<42> net8<43> net8<44> net8<45> net8<46> net8<47> net8<48> 
+ net8<49> net8<50> net8<51> net8<52> net8<53> net8<54> net8<55> net8<56> 
+ net8<57> net8<58> net8<59> net8<60> net8<61> net8<62> net8<63> net035<0> 
+ net035<1> net035<2> net035<3> net035<4> net035<5> net035<6> net035<7> 
+ net035<8> net035<9> net035<10> net035<11> net035<12> net035<13> net035<14> 
+ net035<15> net072<0> net072<1> net072<2> net072<3> net072<4> net072<5> 
+ net072<6> net072<7> net072<8> net072<9> net072<10> net072<11> net072<12> 
+ net072<13> net072<14> net072<15> net072<16> net072<17> net072<18> net072<19> 
+ net072<20> net072<21> net072<22> net072<23> net072<24> net072<25> net072<26> 
+ net072<27> net072<28> net072<29> net072<30> net072<31> net013<0> net013<1> 
+ net013<2> net013<3> net011<0> net011<1> net011<2> net011<3> net011<4> 
+ net011<5> net011<6> net011<7> net011<8> net011<9> net011<10> net011<11> 
+ net011<12> net011<13> net011<14> net011<15> net6<0> net6<1> net6<2> net6<3> 
+ net6<4> net6<5> net6<6> net6<7> net6<8> net6<9> net6<10> net6<11> net6<12> 
+ net6<13> net6<14> net6<15> net6<16> net6<17> net6<18> net6<19> net6<20> 
+ net6<21> net6<22> net6<23> net6<24> net6<25> net6<26> net6<27> net6<28> 
+ net6<29> net6<30> net6<31> net6<32> net6<33> net6<34> net6<35> net6<36> 
+ net6<37> net6<38> net6<39> net6<40> net6<41> net6<42> net6<43> net6<44> 
+ net6<45> net6<46> net6<47> net6<48> net6<49> net6<50> net6<51> net6<52> 
+ net6<53> net6<54> net6<55> net6<56> net6<57> net6<58> net6<59> net6<60> 
+ net6<61> net6<62> net6<63> net036<0> net036<1> net036<2> net036<3> net036<4> 
+ net036<5> net036<6> net036<7> net036<8> net036<9> net036<10> net036<11> 
+ net036<12> net036<13> net036<14> net036<15> vdd vss net014 net09 / 
+ Writedriver
XI3 net027<0> net027<1> net026<0> net026<1> net026<2> net026<3> net026<4> 
+ net026<5> net026<6> net013<0> net013<1> net013<2> net013<3> net025 net024 
+ net10<0> net10<1> net10<2> net10<3> net10<4> net10<5> net10<6> net10<7> 
+ net9<0> net9<1> net9<2> net9<3> net9<4> net9<5> net9<6> net9<7> net9<8> 
+ net9<9> net9<10> net9<11> net9<12> net9<13> net9<14> net9<15> vdd vss net014 
+ net09 / access_decoder
XI4 a<0> a<1> a<2> a<3> a<4> a<5> a<6> a<7> a<8> net027<0> net027<1> net028<0> 
+ net028<1> net028<2> net028<3> net028<4> net090<0> net090<1> net090<2> 
+ net090<3> net026<0> net026<1> net026<2> net026<3> net026<4> net026<5> 
+ net026<6> clk net048 net049 comp net025 net024 net029 net038 net030 inbit 
+ model net078 read set net052 net053 net034 net033 net032 net031 vdd vss wait_ 
+ wrt net014 wrtbuf net09 / master
XI5 net035<0> net035<1> net035<2> net035<3> net035<4> net035<5> net035<6> 
+ net035<7> net035<8> net035<9> net035<10> net035<11> net035<12> net035<13> 
+ net035<14> net035<15> net020<0> net020<1> net020<2> net020<3> net020<4> 
+ net020<5> net020<6> net020<7> net020<8> net020<9> net020<10> net020<11> 
+ net020<12> net020<13> net020<14> net020<15> net020<16> net020<17> net020<18> 
+ net020<19> net020<20> net020<21> net020<22> net020<23> net020<24> net020<25> 
+ net020<26> net020<27> net020<28> net020<29> net020<30> net020<31> net020<32> 
+ net020<33> net020<34> net020<35> net020<36> net020<37> net020<38> net020<39> 
+ net020<40> net020<41> net020<42> net020<43> net020<44> net020<45> net020<46> 
+ net020<47> net020<48> net020<49> net020<50> net020<51> net020<52> net020<53> 
+ net020<54> net020<55> net020<56> net020<57> net020<58> net020<59> net020<60> 
+ net020<61> net020<62> net020<63> net020<64> net020<65> net020<66> net020<67> 
+ net020<68> net020<69> net020<70> net020<71> net020<72> net020<73> net020<74> 
+ net020<75> net020<76> net020<77> net020<78> net020<79> net020<80> net020<81> 
+ net020<82> net020<83> net020<84> net020<85> net020<86> net020<87> net020<88> 
+ net020<89> net020<90> net020<91> net020<92> net020<93> net020<94> net020<95> 
+ net020<96> net020<97> net020<98> net020<99> net020<100> net020<101> 
+ net020<102> net020<103> net020<104> net020<105> net020<106> net020<107> 
+ net020<108> net020<109> net020<110> net020<111> net020<112> net020<113> 
+ net020<114> net020<115> net020<116> net020<117> net020<118> net020<119> 
+ net020<120> net020<121> net020<122> net020<123> net020<124> net020<125> 
+ net020<126> net020<127> net019<0> net019<1> net019<2> net019<3> net019<4> 
+ net019<5> net019<6> net019<7> net019<8> net019<9> net019<10> net019<11> 
+ net019<12> net019<13> net019<14> net019<15> net019<16> net019<17> net019<18> 
+ net019<19> net019<20> net019<21> net019<22> net019<23> net019<24> net019<25> 
+ net019<26> net019<27> net019<28> net019<29> net019<30> net019<31> net019<32> 
+ net019<33> net019<34> net019<35> net019<36> net019<37> net019<38> net019<39> 
+ net019<40> net019<41> net019<42> net019<43> net019<44> net019<45> net019<46> 
+ net019<47> net019<48> net019<49> net019<50> net019<51> net019<52> net019<53> 
+ net019<54> net019<55> net019<56> net019<57> net019<58> net019<59> net019<60> 
+ net019<61> net019<62> net019<63> net019<64> net019<65> net019<66> net019<67> 
+ net019<68> net019<69> net019<70> net019<71> net019<72> net019<73> net019<74> 
+ net019<75> net019<76> net019<77> net019<78> net019<79> net019<80> net019<81> 
+ net019<82> net019<83> net019<84> net019<85> net019<86> net019<87> net019<88> 
+ net019<89> net019<90> net019<91> net019<92> net019<93> net019<94> net019<95> 
+ net019<96> net019<97> net019<98> net019<99> net019<100> net019<101> 
+ net019<102> net019<103> net019<104> net019<105> net019<106> net019<107> 
+ net019<108> net019<109> net019<110> net019<111> net019<112> net019<113> 
+ net019<114> net019<115> net019<116> net019<117> net019<118> net019<119> 
+ net019<120> net019<121> net019<122> net019<123> net019<124> net019<125> 
+ net019<126> net019<127> net015<0> net015<1> net015<2> net015<3> net015<4> 
+ net015<5> net015<6> net015<7> net015<8> net015<9> net015<10> net015<11> 
+ net015<12> net015<13> net015<14> net015<15> net015<16> net015<17> net015<18> 
+ net015<19> net015<20> net015<21> net015<22> net015<23> net015<24> net015<25> 
+ net015<26> net015<27> net015<28> net015<29> net015<30> net015<31> net015<32> 
+ net015<33> net015<34> net015<35> net015<36> net015<37> net015<38> net015<39> 
+ net015<40> net015<41> net015<42> net015<43> net015<44> net015<45> net015<46> 
+ net015<47> net015<48> net015<49> net015<50> net015<51> net015<52> net015<53> 
+ net015<54> net015<55> net015<56> net015<57> net015<58> net015<59> net015<60> 
+ net015<61> net015<62> net015<63> net015<64> net015<65> net015<66> net015<67> 
+ net015<68> net015<69> net015<70> net015<71> net015<72> net015<73> net015<74> 
+ net015<75> net015<76> net015<77> net015<78> net015<79> net015<80> net015<81> 
+ net015<82> net015<83> net015<84> net015<85> net015<86> net015<87> net015<88> 
+ net015<89> net015<90> net015<91> net015<92> net015<93> net015<94> net015<95> 
+ net015<96> net015<97> net015<98> net015<99> net015<100> net015<101> 
+ net015<102> net015<103> net015<104> net015<105> net015<106> net015<107> 
+ net015<108> net015<109> net015<110> net015<111> net015<112> net015<113> 
+ net015<114> net015<115> net015<116> net015<117> net015<118> net015<119> 
+ net015<120> net015<121> net015<122> net015<123> net015<124> net015<125> 
+ net015<126> net015<127> net075<0> net075<1> net075<2> net075<3> net075<4> 
+ net075<5> net075<6> net075<7> net075<8> net075<9> net075<10> net075<11> 
+ net075<12> net075<13> net075<14> net075<15> net075<16> net075<17> net075<18> 
+ net075<19> net075<20> net075<21> net075<22> net075<23> net075<24> net075<25> 
+ net075<26> net075<27> net075<28> net075<29> net075<30> net075<31> net075<32> 
+ net075<33> net075<34> net075<35> net075<36> net075<37> net075<38> net075<39> 
+ net075<40> net075<41> net075<42> net075<43> net075<44> net075<45> net075<46> 
+ net075<47> net075<48> net075<49> net075<50> net075<51> net075<52> net075<53> 
+ net075<54> net075<55> net075<56> net075<57> net075<58> net075<59> net075<60> 
+ net075<61> net075<62> net075<63> net075<64> net075<65> net075<66> net075<67> 
+ net075<68> net075<69> net075<70> net075<71> net075<72> net075<73> net075<74> 
+ net075<75> net075<76> net075<77> net075<78> net075<79> net075<80> net075<81> 
+ net075<82> net075<83> net075<84> net075<85> net075<86> net075<87> net075<88> 
+ net075<89> net075<90> net075<91> net075<92> net075<93> net075<94> net075<95> 
+ net075<96> net075<97> net075<98> net075<99> net075<100> net075<101> 
+ net075<102> net075<103> net075<104> net075<105> net075<106> net075<107> 
+ net075<108> net075<109> net075<110> net075<111> net075<112> net075<113> 
+ net075<114> net075<115> net075<116> net075<117> net075<118> net075<119> 
+ net075<120> net075<121> net075<122> net075<123> net075<124> net075<125> 
+ net075<126> net075<127> net036<0> net036<1> net036<2> net036<3> net036<4> 
+ net036<5> net036<6> net036<7> net036<8> net036<9> net036<10> net036<11> 
+ net036<12> net036<13> net036<14> net036<15> vdd vss net037<0> net037<1> 
+ net037<2> net037<3> net037<4> net037<5> net037<6> net037<7> net037<8> 
+ net037<9> net037<10> net037<11> net037<12> net037<13> net037<14> net037<15> 
+ net037<16> net037<17> net037<18> net037<19> net037<20> net037<21> net037<22> 
+ net037<23> net037<24> net037<25> net037<26> net037<27> net037<28> net037<29> 
+ net037<30> net037<31> / inputbuffer
XI6 net028<0> net028<1> net028<2> net028<3> net028<4> net029 net037<0> 
+ net037<1> net037<2> net037<3> net037<4> net037<5> net037<6> net037<7> 
+ net037<8> net037<9> net037<10> net037<11> net037<12> net037<13> net037<14> 
+ net037<15> net037<16> net037<17> net037<18> net037<19> net037<20> net037<21> 
+ net037<22> net037<23> net037<24> net037<25> net037<26> net037<27> net037<28> 
+ net037<29> net037<30> net037<31> vdd vss / inbuf_decoder
XI7 net035<0> net035<1> net035<2> net035<3> net035<4> net035<5> net035<6> 
+ net035<7> net035<8> net035<9> net035<10> net035<11> net035<12> net035<13> 
+ net035<14> net035<15> net030 net4<0> net4<1> net4<2> net4<3> net4<4> net4<5> 
+ net4<6> net4<7> net4<8> net4<9> net4<10> net4<11> net4<12> net4<13> net4<14> 
+ net4<15> net4<16> net4<17> net4<18> net4<19> net4<20> net4<21> net4<22> 
+ net4<23> net4<24> net4<25> net4<26> net4<27> net4<28> net4<29> net4<30> 
+ net4<31> net4<32> net4<33> net4<34> net4<35> net4<36> net4<37> net4<38> 
+ net4<39> net4<40> net4<41> net4<42> net4<43> net4<44> net4<45> net4<46> 
+ net4<47> net4<48> net4<49> net4<50> net4<51> net4<52> net4<53> net4<54> 
+ net4<55> net4<56> net4<57> net4<58> net4<59> net4<60> net4<61> net4<62> 
+ net4<63> net4<64> net4<65> net4<66> net4<67> net4<68> net4<69> net4<70> 
+ net4<71> net4<72> net4<73> net4<74> net4<75> net4<76> net4<77> net4<78> 
+ net4<79> net4<80> net4<81> net4<82> net4<83> net4<84> net4<85> net4<86> 
+ net4<87> net4<88> net4<89> net4<90> net4<91> net4<92> net4<93> net4<94> 
+ net4<95> net4<96> net4<97> net4<98> net4<99> net4<100> net4<101> net4<102> 
+ net4<103> net4<104> net4<105> net4<106> net4<107> net4<108> net4<109> 
+ net4<110> net4<111> net4<112> net4<113> net4<114> net4<115> net4<116> 
+ net4<117> net4<118> net4<119> net4<120> net4<121> net4<122> net4<123> 
+ net4<124> net4<125> net4<126> net4<127> net5<0> net5<1> net5<2> net5<3> 
+ net5<4> net5<5> net5<6> net5<7> net5<8> net5<9> net5<10> net5<11> net5<12> 
+ net5<13> net5<14> net5<15> net5<16> net5<17> net5<18> net5<19> net5<20> 
+ net5<21> net5<22> net5<23> net5<24> net5<25> net5<26> net5<27> net5<28> 
+ net5<29> net5<30> net5<31> net5<32> net5<33> net5<34> net5<35> net5<36> 
+ net5<37> net5<38> net5<39> net5<40> net5<41> net5<42> net5<43> net5<44> 
+ net5<45> net5<46> net5<47> net5<48> net5<49> net5<50> net5<51> net5<52> 
+ net5<53> net5<54> net5<55> net5<56> net5<57> net5<58> net5<59> net5<60> 
+ net5<61> net5<62> net5<63> net5<64> net5<65> net5<66> net5<67> net5<68> 
+ net5<69> net5<70> net5<71> net5<72> net5<73> net5<74> net5<75> net5<76> 
+ net5<77> net5<78> net5<79> net5<80> net5<81> net5<82> net5<83> net5<84> 
+ net5<85> net5<86> net5<87> net5<88> net5<89> net5<90> net5<91> net5<92> 
+ net5<93> net5<94> net5<95> net5<96> net5<97> net5<98> net5<99> net5<100> 
+ net5<101> net5<102> net5<103> net5<104> net5<105> net5<106> net5<107> 
+ net5<108> net5<109> net5<110> net5<111> net5<112> net5<113> net5<114> 
+ net5<115> net5<116> net5<117> net5<118> net5<119> net5<120> net5<121> 
+ net5<122> net5<123> net5<124> net5<125> net5<126> net5<127> net020<0> 
+ net020<1> net020<2> net020<3> net020<4> net020<5> net020<6> net020<7> 
+ net020<8> net020<9> net020<10> net020<11> net020<12> net020<13> net020<14> 
+ net020<15> net020<16> net020<17> net020<18> net020<19> net020<20> net020<21> 
+ net020<22> net020<23> net020<24> net020<25> net020<26> net020<27> net020<28> 
+ net020<29> net020<30> net020<31> net020<32> net020<33> net020<34> net020<35> 
+ net020<36> net020<37> net020<38> net020<39> net020<40> net020<41> net020<42> 
+ net020<43> net020<44> net020<45> net020<46> net020<47> net020<48> net020<49> 
+ net020<50> net020<51> net020<52> net020<53> net020<54> net020<55> net020<56> 
+ net020<57> net020<58> net020<59> net020<60> net020<61> net020<62> net020<63> 
+ net020<64> net020<65> net020<66> net020<67> net020<68> net020<69> net020<70> 
+ net020<71> net020<72> net020<73> net020<74> net020<75> net020<76> net020<77> 
+ net020<78> net020<79> net020<80> net020<81> net020<82> net020<83> net020<84> 
+ net020<85> net020<86> net020<87> net020<88> net020<89> net020<90> net020<91> 
+ net020<92> net020<93> net020<94> net020<95> net020<96> net020<97> net020<98> 
+ net020<99> net020<100> net020<101> net020<102> net020<103> net020<104> 
+ net020<105> net020<106> net020<107> net020<108> net020<109> net020<110> 
+ net020<111> net020<112> net020<113> net020<114> net020<115> net020<116> 
+ net020<117> net020<118> net020<119> net020<120> net020<121> net020<122> 
+ net020<123> net020<124> net020<125> net020<126> net020<127> net019<0> 
+ net019<1> net019<2> net019<3> net019<4> net019<5> net019<6> net019<7> 
+ net019<8> net019<9> net019<10> net019<11> net019<12> net019<13> net019<14> 
+ net019<15> net019<16> net019<17> net019<18> net019<19> net019<20> net019<21> 
+ net019<22> net019<23> net019<24> net019<25> net019<26> net019<27> net019<28> 
+ net019<29> net019<30> net019<31> net019<32> net019<33> net019<34> net019<35> 
+ net019<36> net019<37> net019<38> net019<39> net019<40> net019<41> net019<42> 
+ net019<43> net019<44> net019<45> net019<46> net019<47> net019<48> net019<49> 
+ net019<50> net019<51> net019<52> net019<53> net019<54> net019<55> net019<56> 
+ net019<57> net019<58> net019<59> net019<60> net019<61> net019<62> net019<63> 
+ net019<64> net019<65> net019<66> net019<67> net019<68> net019<69> net019<70> 
+ net019<71> net019<72> net019<73> net019<74> net019<75> net019<76> net019<77> 
+ net019<78> net019<79> net019<80> net019<81> net019<82> net019<83> net019<84> 
+ net019<85> net019<86> net019<87> net019<88> net019<89> net019<90> net019<91> 
+ net019<92> net019<93> net019<94> net019<95> net019<96> net019<97> net019<98> 
+ net019<99> net019<100> net019<101> net019<102> net019<103> net019<104> 
+ net019<105> net019<106> net019<107> net019<108> net019<109> net019<110> 
+ net019<111> net019<112> net019<113> net019<114> net019<115> net019<116> 
+ net019<117> net019<118> net019<119> net019<120> net019<121> net019<122> 
+ net019<123> net019<124> net019<125> net019<126> net019<127> net015<0> 
+ net015<1> net015<2> net015<3> net015<4> net015<5> net015<6> net015<7> 
+ net015<8> net015<9> net015<10> net015<11> net015<12> net015<13> net015<14> 
+ net015<15> net015<16> net015<17> net015<18> net015<19> net015<20> net015<21> 
+ net015<22> net015<23> net015<24> net015<25> net015<26> net015<27> net015<28> 
+ net015<29> net015<30> net015<31> net015<32> net015<33> net015<34> net015<35> 
+ net015<36> net015<37> net015<38> net015<39> net015<40> net015<41> net015<42> 
+ net015<43> net015<44> net015<45> net015<46> net015<47> net015<48> net015<49> 
+ net015<50> net015<51> net015<52> net015<53> net015<54> net015<55> net015<56> 
+ net015<57> net015<58> net015<59> net015<60> net015<61> net015<62> net015<63> 
+ net015<64> net015<65> net015<66> net015<67> net015<68> net015<69> net015<70> 
+ net015<71> net015<72> net015<73> net015<74> net015<75> net015<76> net015<77> 
+ net015<78> net015<79> net015<80> net015<81> net015<82> net015<83> net015<84> 
+ net015<85> net015<86> net015<87> net015<88> net015<89> net015<90> net015<91> 
+ net015<92> net015<93> net015<94> net015<95> net015<96> net015<97> net015<98> 
+ net015<99> net015<100> net015<101> net015<102> net015<103> net015<104> 
+ net015<105> net015<106> net015<107> net015<108> net015<109> net015<110> 
+ net015<111> net015<112> net015<113> net015<114> net015<115> net015<116> 
+ net015<117> net015<118> net015<119> net015<120> net015<121> net015<122> 
+ net015<123> net015<124> net015<125> net015<126> net015<127> net075<0> 
+ net075<1> net075<2> net075<3> net075<4> net075<5> net075<6> net075<7> 
+ net075<8> net075<9> net075<10> net075<11> net075<12> net075<13> net075<14> 
+ net075<15> net075<16> net075<17> net075<18> net075<19> net075<20> net075<21> 
+ net075<22> net075<23> net075<24> net075<25> net075<26> net075<27> net075<28> 
+ net075<29> net075<30> net075<31> net075<32> net075<33> net075<34> net075<35> 
+ net075<36> net075<37> net075<38> net075<39> net075<40> net075<41> net075<42> 
+ net075<43> net075<44> net075<45> net075<46> net075<47> net075<48> net075<49> 
+ net075<50> net075<51> net075<52> net075<53> net075<54> net075<55> net075<56> 
+ net075<57> net075<58> net075<59> net075<60> net075<61> net075<62> net075<63> 
+ net075<64> net075<65> net075<66> net075<67> net075<68> net075<69> net075<70> 
+ net075<71> net075<72> net075<73> net075<74> net075<75> net075<76> net075<77> 
+ net075<78> net075<79> net075<80> net075<81> net075<82> net075<83> net075<84> 
+ net075<85> net075<86> net075<87> net075<88> net075<89> net075<90> net075<91> 
+ net075<92> net075<93> net075<94> net075<95> net075<96> net075<97> net075<98> 
+ net075<99> net075<100> net075<101> net075<102> net075<103> net075<104> 
+ net075<105> net075<106> net075<107> net075<108> net075<109> net075<110> 
+ net075<111> net075<112> net075<113> net075<114> net075<115> net075<116> 
+ net075<117> net075<118> net075<119> net075<120> net075<121> net075<122> 
+ net075<123> net075<124> net075<125> net075<126> net075<127> net036<0> 
+ net036<1> net036<2> net036<3> net036<4> net036<5> net036<6> net036<7> 
+ net036<8> net036<9> net036<10> net036<11> net036<12> net036<13> net036<14> 
+ net036<15> net034 net033 net032 net031 vdd vss / timegenerate
XI8 net090<0> net090<1> net090<2> net090<3> net040<0> net040<1> net040<2> 
+ net040<3> net040<4> net040<5> net040<6> net040<7> net040<8> net040<9> 
+ net040<10> net040<11> net040<12> net040<13> net040<14> net040<15> net040<16> 
+ net040<17> net040<18> net040<19> net040<20> net040<21> net040<22> net040<23> 
+ net040<24> net040<25> net040<26> net040<27> net040<28> net040<29> net040<30> 
+ net040<31> net011<0> net011<1> net011<2> net011<3> net011<4> net011<5> 
+ net011<6> net011<7> net011<8> net011<9> net011<10> net011<11> net011<12> 
+ net011<13> net011<14> net011<15> net038 net063<0> net063<1> net063<2> 
+ net063<3> net063<4> net063<5> net063<6> net063<7> net063<8> net063<9> 
+ net063<10> net063<11> net063<12> net063<13> net063<14> net063<15> net052 vdd 
+ vss / counter
XI9 net048 net049 d<0> d<1> d<2> d<3> d<4> d<5> d<6> d<7> d<8> d<9> d<10> 
+ d<11> d<12> d<13> d<14> d<15> net011<0> net011<1> net011<2> net011<3> 
+ net011<4> net011<5> net011<6> net011<7> net011<8> net011<9> net011<10> 
+ net011<11> net011<12> net011<13> net011<14> net011<15> net063<0> net063<1> 
+ net063<2> net063<3> net063<4> net063<5> net063<6> net063<7> net063<8> 
+ net063<9> net063<10> net063<11> net063<12> net063<13> net063<14> net063<15> 
+ q<0> q<1> q<2> q<3> q<4> q<5> q<6> q<7> q<8> q<9> q<10> q<11> q<12> q<13> 
+ q<14> q<15> vdd vss / IO
XI11 net040<0> net040<1> net040<2> net040<3> net040<4> net040<5> net040<6> 
+ net040<7> net040<8> net040<9> net040<10> net040<11> net040<12> net040<13> 
+ net040<14> net040<15> net040<16> net040<17> net040<18> net040<19> net040<20> 
+ net040<21> net040<22> net040<23> net040<24> net040<25> net040<26> net040<27> 
+ net040<28> net040<29> net040<30> net040<31> net072<0> net072<1> net072<2> 
+ net072<3> net072<4> net072<5> net072<6> net072<7> net072<8> net072<9> 
+ net072<10> net072<11> net072<12> net072<13> net072<14> net072<15> net072<16> 
+ net072<17> net072<18> net072<19> net072<20> net072<21> net072<22> net072<23> 
+ net072<24> net072<25> net072<26> net072<27> net072<28> net072<29> net072<30> 
+ net072<31> net011<0> net011<1> net011<2> net011<3> net011<4> net011<5> 
+ net011<6> net011<7> net011<8> net011<9> net011<10> net011<11> net011<12> 
+ net011<13> net011<14> net011<15> net078 net052 net053 vdd vss / ADC
.ENDS

.global vdd vss
v_vss vss 0 0
vsu vdd vss 1.2
*.print v(*)

.end