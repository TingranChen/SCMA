// *Spectre Model Format
simulator lang=spectre  insensitive=yes
// * 
// *  no part of this file can be released without the consent of smic.
// *
// ******************************************************************************************
// *         smic 0.18um mixed signal 1p6m 1.8v/3.3v spice model (for hspice only)          *
// ******************************************************************************************
// *
// *  release version    : 1.0
// *
// *  release date       : 04/24/2015
// *
// *  simulation tool    : synopsys star-hspice version c-2010.03
// * 
// *  the valid temperature range is from -40c to 125c
// * model type         :
// *   mosfet           : hspice level 54(bsim4)
// * 
// * simple model name         :
// *        *------------------------------------------------------------*
// *        |     mosfet type    |       1.8v        |        3.3v       |
// *        |============================================================|
// *        |      nmos          | n18_ckt_rf        | n33_ckt_rf        |
// *        *------------------------------------------------------------|
// *        |      pmos          | p18_ckt_rf        | p33_ckt_rf        |
// *        *------------------------------------------------------------|
// *        |      nmos          | dnw18_ckt_rf      | dnw33_ckt_rf      |
// *        *------------------------------------------------------------*
// *        |      pmos          | p18_5t_ckt_rf     | p33_5t_ckt_rf     |
// *        *------------------------------------------------------------*
// *        |      nmos          | dnw18_6t_ckt_rf   | dnw33_6t_ckt_rf   |
// *        *------------------------------------------------------------*
// *
// *    valid temperature range is from -40c to 125c
// *
* 1.8v nmos 
* 1=drain,2=gate,3=source,4=bulk
inline subckt n18_ckt_rf_r (1 2 3 4)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 
**********************************************
+kcgdl=0.5749*Log(lrr*1e6)+1.9162
+kdlc= 0.6197*pwr(lrr*1e6,-0.336)
+Cgd_rf = max((0.1754*pwr(lrr*1000000,0.8196)*wrr*1000000+0.2349*pwr(lrr*1000000,2.0815)+0.35)*nfr*1e-15*(0.4736*pwr(nfr,-1.785)+0.999),1e-18)  
+Cgs_rf = max((0.0312*exp(-2.228*lrr*1e6)*wrr*1e6+0.1664*log(lrr*1e6)+0.6883)*nfr*1e-15*(2.3304*pwr(nfr,-0.836)+0.88),1e-18)
+Cds_rf = max(max((-0.192*Log(lrr*1e6)-0.1941)*wrr*1e6+1/(0.00000264*pwr(lrr*1e6,-7.76)+10.92),0.03)*nfr*1e-15,1e-18)
+Rg_rf =  max(1/(0.0327*pwr(lrr*1000000,1.0167)*pwr(wrr*1000000,0.3525*EXP(1.1485*lrr*1000000))*(nfr+3)),1e-3) 
+Rsub1_rf = max((-3.6736*nfr+179.52)*(1/(27.288*pwr(lrr*1e6,3.3796)+0.75)),5)
+Rsub2_rf = 35
+Djdb_AREA_rf = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf   = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*11.6749)                                                                                          
+Djsb_AREA_rf = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf   = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*11.6749)  
**********************************************
Lgate       ( 2 20) inductor  l=1p                        m=mrr
Rgate       (20 21) resistor  r=Rg_rf*(1+drg_n18_rf)      m=mrr
Cgd_ext     (21 11) capacitor c=Cgd_rf*(1+dcgdext_n18_rf) m=mrr
Cgs_ext     (21 31) capacitor c=Cgs_rf*(1+dcgsext_n18_rf) m=mrr
Cds_ext     (15 31) capacitor c=Cds_rf                    m=mrr
Rds         (11 15) resistor  r=10                        m=mrr
Ldrain       (1 11) inductor  l=1p                        m=mrr
Lsource      (3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (12 11) ndio18_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (32 31) ndio18_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
**********************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
**********************************************
n18_ckt_rf_r (11 21 31 41) n18_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model n18_ckt_r bsim4 type = n
**********************************************************************************************                                                                            
*                              1.8V CORE NMOS MODEL                               *                                                                            
**********************************************************************************************                                                                            
*                                                                                                                                            
*                                                                                                                                                              
* GENERAL PARAMETERS                                                                                                                                           
*                                                                                                                                                              
***************************************************************************                                                                                    
*             Model Selector Parameter                                                                                                                         
***************************************************************************                                                                                    
+level        = 54                version      = 4.5               binunit      = 2                                                                            
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                                                                            
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                                                                            
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                                                                            
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                                                                            
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                                                                            
+igcmod       = 1                 igbmod       = 1                 wpemod       = 0                                                                            
                                                                                                                                                               
***************************************************************************                                                                                    
*             Geometry Range Parameter                                                                                                                         
***************************************************************************                                                                                    
+lmin         = 1.5e-007          lmax         = 0.0001            wmin         = 1.9e-007          
+wmax         = 0.0001
***************************************************************************                                                                                    
*             Process Parameter                                                                                                                                
***************************************************************************                                                                                    
+epsrox       = 3.9                                                                                                                                            
+toxe         = 4.19e-009+dtoxe_n18_rf_mismatch                                                                                                                        
+dtox         = 3.36e-010         xj           = 1.6e-007          ndep         = 1.4563e+017                                                                  
+ngate        = 3e+020            nsd          = 1e+020            rsh          = 7.6
***************************************************************************                                                                                    
*             dW and dL Parameter                                                                                                                              
***************************************************************************                                                                                    
+wl           = 0                 wln          = 1                 ww           = -2.7e-015         
+wwn          = 1                 wwl          = -8e-022           ll           = -7e-016           
+lln          = 1                 lw           = -3.5e-015         lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 wint         = 1.6229e-008       lint         = 9e-009 
***************************************************************************                                                                                    
*             Layout-Dependent Parasitics Model Parameter                                                                                                      
***************************************************************************                                                                                    
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                                                                            
+xgw          =0.31e-6            xgl          =-1.6e-008          ngcon        =2       
+xl           = -1.6e-008+dxl_n18_rf                                                                                                                         
+xw           = 4.2e-008+dxw_n18_rf
***************************************************************************                                                                                    
*             BASIC: Vth Related  Parameter                                                                                                                    
***************************************************************************                                                                                          
+vth0         = 0.4185+dvth0_n18_rf_mismatch                                                             
+lvth0        = -1.495e-008+dlvth0_n18_rf                                                       
+wvth0        = -1.16e-008+dwvth0_n18_rf                                                        
+pvth0        = 1.8e-015+dpvth0_n18_rf                                                          
+vfb          = -1                phin         = 0.077042          k1           = 0.57819           
+wk1          = -1.7e-008         k2           = 0.0024336         lk2          = -1e-009           
+wk2          = 2e-009            pk2          = 1.4699e-015       k3           = 3                 
+k3b          = 3.76              w0           = 1.5e-006          lpe0         = 1.8e-007          
+llpe0        = 1.1e-016          lpeb         = 0                 vbm          = -3                
+dvt0         = 1.14              ldvt0        = -6.124e-008       dvt1         = 0.22              
+ldvt1        = 2e-009            dvt2         = -0.02944          dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            dwg          = 0                 dwb          = 0
***************************************************************************                                                                                    
*             BASIC: Mobility Related Parameter                                                                                                                
***************************************************************************                                                                                    
+u0           = 0.028012+du0_n18_rf_mismatch                                                            
+lu0          = 5.4e-010+dlu0_n18_rf                                                           
+wu0          = -4.51e-010+dwu0_n18_rf                                                         
+pu0          = 4.6575e-016+dpu0_n18_rf                                                        
+ua           = -1.8869e-009      lua          = -3e-017           wua          = 7.6568e-017       
+pua          = 6.4915e-024       ub           = 3.515e-018        lub          = 2.92e-026         
+wub          = -1.274e-025       pub          = -7.86e-033        uc           = 1.4426e-010       
+luc          = 2.1688e-018       wuc          = -1.2768e-017      puc          = 8e-025            
+ud           = 0                 eu           = 1.67              
+vsat         = 70000+dvsat_n18_rf_mismatch                                                             
+lvsat        = 0.0006+dlvsat_n18_rf                                                           
+pvsat        = 5.2036e-010+dpvsat_n18_rf                                                      
+a0           = 1.6               la0          = -4e-007           pa0          = 5e-014            
+ags          = 0.56              lags         = 1.5e-007          wags         = -3e-008           
+pags         = 6e-014            b0           = 0                 b1           = 0                 
+keta         = -0.045548         lketa        = -7.6454e-009      wketa        = 1.0136e-008       
+pketa        = -1e-015           a1           = 0                 a2           = 0.99                                                                         
***************************************************************************  
*             BASIC: Subthreshold Related Parameter                           
***************************************************************************    
+voff         = -0.15+dvoff_n18_rf                                                             
+pvoff        = -5e-016           voffl        = 0                 minv         = 0                 
+nfactor      = 1                 eta0         = 0.14              peta0        = -6e-016           
+etab         = -0.07             petab        = 3.6e-015          dsub         = 0.56              
+cit          = 0.00065           lcit         = 1.6e-010          pcit         = -1e-018           
+cdsc         = 0                 cdscb        = 0                 cdscd        = 0.0001
***************************************************************************                                                                                    
*             BASIC: Output Resistance Related Parameter                                                                                                       
***************************************************************************                                                                                    
+pclm         = 0.31747           ppclm        = 4e-015            pdiblc1      = 0.04              
+pdiblc2      = 0.002             pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 3.45e+008         pscbe2       = 1e-006            pvag         = 0                 
+delta        = 0.001             pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 lambda       = 0 
***************************************************************************                                                                                    
*             Asymmetric and Bias-Dependent                                                                                                                    
***************************************************************************                                                                                    
+rdsw         = 90                rdswmin      = 0                 rdw          = 47                
+rdwmin       = 0                 rsw          = 47                rswmin       = 0                 
+prwg         = 0                 prwb         = 0                 wr           = 1  
***************************************************************************                                                                                    
*             Impact Ionization Current Model Parameters                                                                                                       
***************************************************************************                                                                                    
+alpha0       = 0                 alpha1       = 4.1739            lalpha1      = 2e-007            
+walpha1      = 4.64e-008         palpha1      = 2.5e-014          beta0        = 15.901    
***************************************************************************                                                                                    
*             Gate Dielectric Tunneling Current                                                                                                                
***************************************************************************                                                                                    
+aigbacc      = 0.43              bigbacc      = 0.054             cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0088021         bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.015123          bigc         = 0.0017647         cigc         = 0.0702            
+dlcig        = 1e-012            aigsd        = 0.0038304         waigsd       = -2e-010           
+paigsd       = -5e-018           bigsd        = 0.00030435        cigsd        = 0.19301           
+nigc         = 1.288             poxedge      = 1                 pigcd        = 1                 
+ntox         = 1                 toxref       = 3e-009          
***************************************************************************                                                                                    
*             GIDL Effect Parameters                                                                                                                           
***************************************************************************                                                                                    
+agidl        = 8.5074e-007       wagidl       = 2e-013            bgidl        = 2.9037e+009       
+wbgidl       = -50               cgidl        = 0.1               egidl        = 0.1        
***************************************************************************                                                                                    
*             Flicker Noise Model Parameter                                                                                                                    
***************************************************************************                                                                                    
+noia         = 6.24173e+041      noib         = 1.42569e+022      noic         = 6.62e+008                                                                    
+em           = 54761.2           ef           = 0.98              lintnoi      = -2e-008                                                                      
+ntnoi        = 1 
***************************************************************************                                                                                    
*             High-Speed RF Model Parameters                                                                                                                   
***************************************************************************                                                                                    
+rnoia=(-2.6579E-01*log(lrr)-3.3425E+00) tnoia=(1.8380E+06*log(lrr)+3.1801E+07) rnoib=0 tnoib=2e6                                                                                                                                                                                                                                    
***************************************************************************                                                                                    
*             Capacitance Parameter                                                                                                                            
***************************************************************************                                                                                    
+xpart        = 0                                                                                                                                              
+cgdo         = 1.8e-010+dcgdo_n18_rf                                                                                                                        
+cgso         = 1.8e-010+dcgdo_n18_rf                                                                                                                        
+cgbo         = 0                                                                                                                                              
+cgdl         = 9e-011*kcgdl+dcgdl_n18_rf                                                                                                                          
+cgsl         = 9e-011*kcgdl+dcgdl_n18_rf                                                                                                                          
+cf           = (8.54e-011+dcf_n18_rf)                                                                                                                         
+clc          = 0                 cle          = 0.6               dlc          = 2.8339e-008*kdlc                                                                  
+dwc          = 0                 vfbcv        = -1                noff         = 1.6804                                                                       
+lnoff        = 1e-007            voffcv       = -0.020304         lvoffcv      = -2.088e-009                                                                  
+acde         = 0.384             moin         = 8                                                                                                       

*+dwc          = 0                 vfbcv        = -1                noff         = 1.6804                                                                     
*+lnoff        = 1e-007            voffcv       = -0.015        lvoffcv      = 0   
*+lnoff        = 1e-007            voffcv       = -0.02        lvoffcv      = 0                                                                
                                                             
*************************************************************************** 
*             Souce|Drain Junction Diode Model Parameter                     
***************************************************************************   
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.5              jss          = 1.1508e-006       jsws         = 1.4205e-014       
+jswgs        = 1.134e-013        jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 2e-008            
+jtsswgd      = 6e-009            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                                                                                                                                               
+cjs          = 0                                                                                                                        
+cjsws        = 0                                                                                                                     
+cjswgs       = 0                                                                                                                    
+mjs          = 0.34744           mjsws        = 0.19672           mjswgs       = 0.84898           
+pbs          = 0.70413           pbsws        = 0.58719           pbswgs       = 1.6255                                                                                                                                                               
***************************************************************************                                                                                    
*             Temperature coefficient                                                                                                                          
***************************************************************************                                                                                    
+tnom         = 25                ute          = -1.4012           lute         = 1.48e-008         
+kt1          = -0.24949          kt1l         = -2.9274e-009      kt2          = -0.05             
+wkt2         = 4e-009            ua1          = 1.76e-009         wua1         = -1.1e-016         
+pua1         = 1.625e-023        ub1          = -1.9392e-018      lub1         = -8.232e-026       
+wub1         = 1e-026            pub1         = -3.12e-033        uc1          = 1.124e-010        
+luc1         = -1.62e-017        puc1         = -3e-024           at           = 31820             
+pat          = -2.1e-010         prt          = 0                 njs          = 1.1294            
+xtis         = 3                 tpb          = 0.001             tpbsw        = 0.000868          
+tpbswg       = 0.0015811         tcj          = 0.00083836        tcjsw        = 0.0014935         
+tcjswg       = 0.0006583         tvoff        = 0                                                                                                               
***************************************************************************                                                                                    
*             Stress Effect Related Parameter                                                                                                                  
***************************************************************************                                                                                    
+saref        = 4.48e-006         sbref        = 4.48e-006         wlod         = 0                 
+ku0          = -4.5e-008         kvsat        = 1                 tku0         = 0                 
+lku0         = 7e-007            wku0         = 5e-007            pku0         = 7e-013            
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 3.5e-009          
+lkvth0       = -6e-008           wkvth0       = 1e-007            pkvth0       = 2e-014            
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                                                                                                                                                                
***************************************************************************                                                                                    
*             Well Proximity Effect Model Parameters                                                                                                           
***************************************************************************                                                                                    
+web          = 0                 wec          = 0                 kvth0we      = 0                                                                            
+k2we         = 0                 ku0we        = 0                 scref        = 1e-006                                                                       
***rf***                                                                                                                                                       
+ XRCRG1  = 12              XRCRG2  = 1                                                                                                                      
+ RSHG    =(rshg_n18_rf)                                                                                                                                               
******************************************************
* **
model ndio18_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 1.1508e-006 isw = 1.4205e-014 vb = 11.5 ibv = 55.6 
+n = 1.1294 ns = 1.1294 rs = 5.0328e-010 
+cj = 0.00098714+dcj_n18_rf cjsw = 5.8272e-011*0.7+dcjsw_n18_rf vj = 0.70413 vjsw = 0.58719 
+fcs = 0 mj = 0.34744 mjsw = 0.2 fc = 0 
+tlev = 1 tlevc = 1 trs = 0.0019296 xti = 3 
+cta = 0.00083836 ctp = 0.001 pta = 0.001395 ptp = 0.000868 
+eg = 1.16  tcv = -0.0004
* *                           

ends n18_ckt_rf_r


* 1.8v nmos in dnw with 4 ports
* 1=drain,2=gate,3=source,4=bulk
inline subckt dnw18_ckt_rf_r (1 2 3 4)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 
**********************************************
+kcgdl=0.5749*Log(lrr*1e6)+1.9162
+kdlc= 0.6197*pwr(lrr*1e6,-0.336)
+Cgd_rf = max((0.1754*pwr(lrr*1000000,0.8196)*wrr*1000000+0.2349*pwr(lrr*1000000,2.0815)+0.35)*nfr*1e-15*(0.4736*pwr(nfr,-1.785)+0.999),1e-18)  
+Cgs_rf = max((0.0312*exp(-2.228*lrr*1e6)*wrr*1e6+0.1664*log(lrr*1e6)+0.6883)*nfr*1e-15*(2.3304*pwr(nfr,-0.836)+0.88),1e-18)
+Cds_rf = max(max((-0.192*Log(lrr*1e6)-0.1941)*wrr*1e6+1/(0.00000264*pwr(lrr*1e6,-7.76)+10.92),0.03)*nfr*1e-15,1e-18)
+Rg_rf =  max(1/(0.0327*pwr(lrr*1000000,1.0167)*pwr(wrr*1000000,0.3525*EXP(1.1485*lrr*1000000))*(nfr+3)),1e-3) 
+Rsub1_rf = max((-3.6736*nfr+179.52)*(1/(27.288*pwr(lrr*1e6,3.3796)+0.75)),5)
+Rsub2_rf = 35
+Djdb_AREA_rf = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf   = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*11.6749)                                                                                          
+Djsb_AREA_rf = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf   = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*11.6749)  
**********************************************
Lgate       ( 2 20) inductor  l=1p                        m=mrr
Rgate       (20 21) resistor  r=Rg_rf*(1+drg_n18_rf)      m=mrr
Cgd_ext     (21 11) capacitor c=Cgd_rf*(1+dcgdext_n18_rf) m=mrr
Cgs_ext     (21 31) capacitor c=Cgs_rf*(1+dcgsext_n18_rf) m=mrr
Cds_ext     (15 31) capacitor c=Cds_rf                    m=mrr
Rds         (11 15) resistor  r=10                        m=mrr
Ldrain       (1 11) inductor  l=1p                        m=mrr
Lsource      (3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (12 11) ndio18_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (32 31) ndio18_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
**********************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
**********************************************
dnw18_ckt_rf_r (11 21 31 41) n18_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model n18_ckt_r bsim4 type = n
**********************************************************************************************                                                                            
*                              1.8V CORE NMOS MODEL                               *                                                                            
**********************************************************************************************                                                                            
*                                                                                                                                            
*                                                                                                                                                              
* GENERAL PARAMETERS                                                                                                                                           
*                                                                                                                                                              
***************************************************************************                                                                                    
*             Model Selector Parameter                                                                                                                         
***************************************************************************                                                                                    
+level        = 54                version      = 4.5               binunit      = 2                                                                            
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                                                                            
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                                                                            
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                                                                            
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                                                                            
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                                                                            
+igcmod       = 1                 igbmod       = 1                 wpemod       = 0                                                                            
                                                                                                                                                               
***************************************************************************                                                                                    
*             Geometry Range Parameter                                                                                                                         
***************************************************************************                                                                                    
+lmin         = 1.5e-007          lmax         = 0.0001            wmin         = 1.9e-007          
+wmax         = 0.0001
***************************************************************************                                                                                    
*             Process Parameter                                                                                                                                
***************************************************************************                                                                                    
+epsrox       = 3.9                                                                                                                                            
+toxe         = 4.19e-009+dtoxe_n18_rf_mismatch                                                                                                                        
+dtox         = 3.36e-010         xj           = 1.6e-007          ndep         = 1.4563e+017                                                                  
+ngate        = 3e+020            nsd          = 1e+020            rsh          = 7.6
***************************************************************************                                                                                    
*             dW and dL Parameter                                                                                                                              
***************************************************************************                                                                                    
+wl           = 0                 wln          = 1                 ww           = -2.7e-015         
+wwn          = 1                 wwl          = -8e-022           ll           = -7e-016           
+lln          = 1                 lw           = -3.5e-015         lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 wint         = 1.6229e-008       lint         = 9e-009 
***************************************************************************                                                                                    
*             Layout-Dependent Parasitics Model Parameter                                                                                                      
***************************************************************************                                                                                    
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                                                                            
+xgw          =0.31e-6            xgl          =-1.6e-008          ngcon        =2       
+xl           = -1.6e-008+dxl_n18_rf                                                                                                                         
+xw           = 4.2e-008+dxw_n18_rf
***************************************************************************                                                                                    
*             BASIC: Vth Related  Parameter                                                                                                                    
***************************************************************************                                                                                          
+vth0         = 0.4185+dvth0_n18_rf_mismatch                                                             
+lvth0        = -1.495e-008+dlvth0_n18_rf                                                       
+wvth0        = -1.16e-008+dwvth0_n18_rf                                                        
+pvth0        = 1.8e-015+dpvth0_n18_rf                                                          
+vfb          = -1                phin         = 0.077042          k1           = 0.57819           
+wk1          = -1.7e-008         k2           = 0.0024336         lk2          = -1e-009           
+wk2          = 2e-009            pk2          = 1.4699e-015       k3           = 3                 
+k3b          = 3.76              w0           = 1.5e-006          lpe0         = 1.8e-007          
+llpe0        = 1.1e-016          lpeb         = 0                 vbm          = -3                
+dvt0         = 1.14              ldvt0        = -6.124e-008       dvt1         = 0.22              
+ldvt1        = 2e-009            dvt2         = -0.02944          dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            dwg          = 0                 dwb          = 0
***************************************************************************                                                                                    
*             BASIC: Mobility Related Parameter                                                                                                                
***************************************************************************                                                                                    
+u0           = 0.028012+du0_n18_rf_mismatch                                                            
+lu0          = 5.4e-010+dlu0_n18_rf                                                           
+wu0          = -4.51e-010+dwu0_n18_rf                                                         
+pu0          = 4.6575e-016+dpu0_n18_rf                                                        
+ua           = -1.8869e-009      lua          = -3e-017           wua          = 7.6568e-017       
+pua          = 6.4915e-024       ub           = 3.515e-018        lub          = 2.92e-026         
+wub          = -1.274e-025       pub          = -7.86e-033        uc           = 1.4426e-010       
+luc          = 2.1688e-018       wuc          = -1.2768e-017      puc          = 8e-025            
+ud           = 0                 eu           = 1.67              
+vsat         = 70000+dvsat_n18_rf_mismatch                                                             
+lvsat        = 0.0006+dlvsat_n18_rf                                                           
+pvsat        = 5.2036e-010+dpvsat_n18_rf                                                      
+a0           = 1.6               la0          = -4e-007           pa0          = 5e-014            
+ags          = 0.56              lags         = 1.5e-007          wags         = -3e-008           
+pags         = 6e-014            b0           = 0                 b1           = 0                 
+keta         = -0.045548         lketa        = -7.6454e-009      wketa        = 1.0136e-008       
+pketa        = -1e-015           a1           = 0                 a2           = 0.99                                                                         
***************************************************************************  
*             BASIC: Subthreshold Related Parameter                           
***************************************************************************    
+voff         = -0.15+dvoff_n18_rf                                                             
+pvoff        = -5e-016           voffl        = 0                 minv         = 0                 
+nfactor      = 1                 eta0         = 0.14              peta0        = -6e-016           
+etab         = -0.07             petab        = 3.6e-015          dsub         = 0.56              
+cit          = 0.00065           lcit         = 1.6e-010          pcit         = -1e-018           
+cdsc         = 0                 cdscb        = 0                 cdscd        = 0.0001
***************************************************************************                                                                                    
*             BASIC: Output Resistance Related Parameter                                                                                                       
***************************************************************************                                                                                    
+pclm         = 0.31747           ppclm        = 4e-015            pdiblc1      = 0.04              
+pdiblc2      = 0.002             pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 3.45e+008         pscbe2       = 1e-006            pvag         = 0                 
+delta        = 0.001             pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 lambda       = 0 
***************************************************************************                                                                                    
*             Asymmetric and Bias-Dependent                                                                                                                    
***************************************************************************                                                                                    
+rdsw         = 90                rdswmin      = 0                 rdw          = 47                
+rdwmin       = 0                 rsw          = 47                rswmin       = 0                 
+prwg         = 0                 prwb         = 0                 wr           = 1  
***************************************************************************                                                                                    
*             Impact Ionization Current Model Parameters                                                                                                       
***************************************************************************                                                                                    
+alpha0       = 0                 alpha1       = 4.1739            lalpha1      = 2e-007            
+walpha1      = 4.64e-008         palpha1      = 2.5e-014          beta0        = 15.901    
***************************************************************************                                                                                    
*             Gate Dielectric Tunneling Current                                                                                                                
***************************************************************************                                                                                    
+aigbacc      = 0.43              bigbacc      = 0.054             cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0088021         bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.015123          bigc         = 0.0017647         cigc         = 0.0702            
+dlcig        = 1e-012            aigsd        = 0.0038304         waigsd       = -2e-010           
+paigsd       = -5e-018           bigsd        = 0.00030435        cigsd        = 0.19301           
+nigc         = 1.288             poxedge      = 1                 pigcd        = 1                 
+ntox         = 1                 toxref       = 3e-009          
***************************************************************************                                                                                    
*             GIDL Effect Parameters                                                                                                                           
***************************************************************************                                                                                    
+agidl        = 8.5074e-007       wagidl       = 2e-013            bgidl        = 2.9037e+009       
+wbgidl       = -50               cgidl        = 0.1               egidl        = 0.1        
***************************************************************************                                                                                    
*             Flicker Noise Model Parameter                                                                                                                    
***************************************************************************                                                                                    
+noia         = 6.24173e+041      noib         = 1.42569e+022      noic         = 6.62e+008                                                                    
+em           = 54761.2           ef           = 0.98              lintnoi      = -2e-008                                                                      
+ntnoi        = 1 
***************************************************************************                                                                                    
*             High-Speed RF Model Parameters                                                                                                                   
***************************************************************************                                                                                    
+rnoia=(-2.6579E-01*log(lrr)-3.3425E+00) tnoia=(1.8380E+06*log(lrr)+3.1801E+07) rnoib=0 tnoib=2e6                                                                                                                                                                
***************************************************************************                                                                                    
*             Capacitance Parameter                                                                                                                            
***************************************************************************                                                                                    
+xpart        = 0                                                                                                                                              
+cgdo         = 1.8e-010+dcgdo_n18_rf                                                                                                                        
+cgso         = 1.8e-010+dcgdo_n18_rf                                                                                                                        
+cgbo         = 0                                                                                                                                              
+cgdl         = 9e-011*kcgdl+dcgdl_n18_rf                                                                                                                          
+cgsl         = 9e-011*kcgdl+dcgdl_n18_rf                                                                                                                          
+cf           = (8.54e-011+dcf_n18_rf)                                                                                                                         
+clc          = 0                 cle          = 0.6               dlc          = 2.8339e-008*kdlc                                                                  
+dwc          = 0                 vfbcv        = -1                noff         = 1.6804                                                                       
+lnoff        = 1e-007            voffcv       = -0.020304         lvoffcv      = -2.088e-009                                                                  
+acde         = 0.384             moin         = 8                                                                                                       

*+dwc          = 0                 vfbcv        = -1                noff         = 1.6804                                                                     
*+lnoff        = 1e-007            voffcv       = -0.015        lvoffcv      = 0   
*+lnoff        = 1e-007            voffcv       = -0.02        lvoffcv      = 0                                                                
                                                             
*************************************************************************** 
*             Souce|Drain Junction Diode Model Parameter                     
***************************************************************************   
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.5              jss          = 1.1508e-006       jsws         = 1.4205e-014       
+jswgs        = 1.134e-013        jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 2e-008            
+jtsswgd      = 6e-009            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                                                                                                                                               
+cjs          = 0                                                                                                                        
+cjsws        = 0                                                                                                                     
+cjswgs       = 0                                                                                                                    
+mjs          = 0.34744           mjsws        = 0.19672           mjswgs       = 0.84898           
+pbs          = 0.70413           pbsws        = 0.58719           pbswgs       = 1.6255                                                                                                                                                               
***************************************************************************                                                                                    
*             Temperature coefficient                                                                                                                          
***************************************************************************                                                                                    
+tnom         = 25                ute          = -1.4012           lute         = 1.48e-008         
+kt1          = -0.24949          kt1l         = -2.9274e-009      kt2          = -0.05             
+wkt2         = 4e-009            ua1          = 1.76e-009         wua1         = -1.1e-016         
+pua1         = 1.625e-023        ub1          = -1.9392e-018      lub1         = -8.232e-026       
+wub1         = 1e-026            pub1         = -3.12e-033        uc1          = 1.124e-010        
+luc1         = -1.62e-017        puc1         = -3e-024           at           = 31820             
+pat          = -2.1e-010         prt          = 0                 njs          = 1.1294            
+xtis         = 3                 tpb          = 0.001             tpbsw        = 0.000868          
+tpbswg       = 0.0015811         tcj          = 0.00083836        tcjsw        = 0.0014935         
+tcjswg       = 0.0006583         tvoff        = 0                                                                                                               
***************************************************************************                                                                                    
*             Stress Effect Related Parameter                                                                                                                  
***************************************************************************                                                                                    
+saref        = 4.48e-006         sbref        = 4.48e-006         wlod         = 0                 
+ku0          = -4.5e-008         kvsat        = 1                 tku0         = 0                 
+lku0         = 7e-007            wku0         = 5e-007            pku0         = 7e-013            
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 3.5e-009          
+lkvth0       = -6e-008           wkvth0       = 1e-007            pkvth0       = 2e-014            
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                                                                                                                                                                
***************************************************************************                                                                                    
*             Well Proximity Effect Model Parameters                                                                                                           
***************************************************************************                                                                                    
+web          = 0                 wec          = 0                 kvth0we      = 0                                                                            
+k2we         = 0                 ku0we        = 0                 scref        = 1e-006                                                                       
***rf***                                                                                                                                                       
+ XRCRG1  = 12              XRCRG2  = 1                                                                                                                      
+ RSHG    =(rshg_n18_rf)                                                                                                                                               
******************************************************
* **
model ndio18_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 1.1508e-006 isw = 1.4205e-014 vb = 11.5 ibv = 55.6 
+n = 1.1294 ns = 1.1294 rs = 5.0328e-010 
+cj = 0.00098714+dcj_n18_rf cjsw = 5.8272e-011*0.7+dcjsw_n18_rf vj = 0.70413 vjsw = 0.58719 
+fcs = 0 mj = 0.34744 mjsw = 0.2 fc = 0 
+tlev = 1 tlevc = 1 trs = 0.0019296 xti = 3 
+cta = 0.00083836 ctp = 0.001 pta = 0.001395 ptp = 0.000868 
+eg = 1.16  tcv = -0.0004
* *                           

ends dnw18_ckt_rf_r


* 1.8v nmos in dnw with 6 ports
* 1=drain,2=gate,3=source,4=bulk,5=dnw,6=psub
inline subckt dnw18_6t_ckt_rf_r (1 2 3 4 5 6)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 arpwr=51.8e-12 pjpwr=28.8e-6 ardnwr=77.4e-12 pjdnwr=35.2e-6 
**********************************************
+kcgdl=0.5749*Log(lrr*1e6)+1.9162
+kdlc= 0.6197*pwr(lrr*1e6,-0.336)
+Cgd_rf = max((0.1754*pwr(lrr*1000000,0.8196)*wrr*1000000+0.2349*pwr(lrr*1000000,2.0815)+0.35)*nfr*1e-15*(0.4736*pwr(nfr,-1.785)+0.999),1e-18)  
+Cgs_rf = max((0.0312*exp(-2.228*lrr*1e6)*wrr*1e6+0.1664*log(lrr*1e6)+0.6883)*nfr*1e-15*(2.3304*pwr(nfr,-0.836)+0.88),1e-18)
+Cds_rf = max(max((-0.192*Log(lrr*1e6)-0.1941)*wrr*1e6+1/(0.00000264*pwr(lrr*1e6,-7.76)+10.92),0.03)*nfr*1e-15,1e-18)
+Rg_rf =  max(1/(0.0327*pwr(lrr*1000000,1.0167)*pwr(wrr*1000000,0.3525*EXP(1.1485*lrr*1000000))*(nfr+3)),1e-3) 
+Rsub1_rf = max((-3.6736*nfr+179.52)*(1/(27.288*pwr(lrr*1e6,3.3796)+0.75)),5)
+Rsub2_rf = 35
+Djdb_AREA_rf = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf   = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*11.6749)                                                                                          
+Djsb_AREA_rf = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf   = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*11.6749)  
**********************************************
Lgate       ( 2 20) inductor  l=1p                        m=mrr
Rgate       (20 21) resistor  r=Rg_rf*(1+drg_n18_rf)      m=mrr
Cgd_ext     (21 11) capacitor c=Cgd_rf*(1+dcgdext_n18_rf) m=mrr
Cgs_ext     (21 31) capacitor c=Cgs_rf*(1+dcgsext_n18_rf) m=mrr
Cds_ext     (15 31) capacitor c=Cds_rf                    m=mrr
Rds         (11 15) resistor  r=10                        m=mrr
Ldrain       (1 11) inductor  l=1p                        m=mrr
Lsource      (3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (12 11) ndio18_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (32 31) ndio18_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
djbdn  (4 5) diobpw_rf area=arpwr pj=pjpwr m=mrr
djpsub (6 5) dnwdio_rf area=ardnwr pj=pjdnwr m=mrr
**********************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
**********************************************
dnw18_6t_ckt_rf_r (11 21 31 41) n18_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model n18_ckt_r bsim4 type = n
**********************************************************************************************                                                                            
*                              1.8V CORE NMOS MODEL                               *                                                                            
**********************************************************************************************                                                                            
*                                                                                                                                            
*                                                                                                                                                              
* GENERAL PARAMETERS                                                                                                                                           
*                                                                                                                                                              
***************************************************************************                                                                                    
*             Model Selector Parameter                                                                                                                         
***************************************************************************                                                                                    
+level        = 54                version      = 4.5               binunit      = 2                                                                            
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                                                                            
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                                                                            
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                                                                            
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                                                                            
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                                                                            
+igcmod       = 1                 igbmod       = 1                 wpemod       = 0                                                                            
                                                                                                                                                               
***************************************************************************                                                                                    
*             Geometry Range Parameter                                                                                                                         
***************************************************************************                                                                                    
+lmin         = 1.5e-007          lmax         = 0.0001            wmin         = 1.9e-007          
+wmax         = 0.0001
***************************************************************************                                                                                    
*             Process Parameter                                                                                                                                
***************************************************************************                                                                                    
+epsrox       = 3.9                                                                                                                                            
+toxe         = 4.19e-009+dtoxe_n18_rf_mismatch                                                                                                                        
+dtox         = 3.36e-010         xj           = 1.6e-007          ndep         = 1.4563e+017                                                                  
+ngate        = 3e+020            nsd          = 1e+020            rsh          = 7.6
***************************************************************************                                                                                    
*             dW and dL Parameter                                                                                                                              
***************************************************************************                                                                                    
+wl           = 0                 wln          = 1                 ww           = -2.7e-015         
+wwn          = 1                 wwl          = -8e-022           ll           = -7e-016           
+lln          = 1                 lw           = -3.5e-015         lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 wint         = 1.6229e-008       lint         = 9e-009 
***************************************************************************                                                                                    
*             Layout-Dependent Parasitics Model Parameter                                                                                                      
***************************************************************************                                                                                    
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                                                                            
+xgw          =0.31e-6            xgl          =-1.6e-008          ngcon        =2       
+xl           = -1.6e-008+dxl_n18_rf                                                                                                                         
+xw           = 4.2e-008+dxw_n18_rf
***************************************************************************                                                                                    
*             BASIC: Vth Related  Parameter                                                                                                                    
***************************************************************************                                                                                          
+vth0         = 0.4185+dvth0_n18_rf_mismatch                                                             
+lvth0        = -1.495e-008+dlvth0_n18_rf                                                       
+wvth0        = -1.16e-008+dwvth0_n18_rf                                                        
+pvth0        = 1.8e-015+dpvth0_n18_rf                                                          
+vfb          = -1                phin         = 0.077042          k1           = 0.57819           
+wk1          = -1.7e-008         k2           = 0.0024336         lk2          = -1e-009           
+wk2          = 2e-009            pk2          = 1.4699e-015       k3           = 3                 
+k3b          = 3.76              w0           = 1.5e-006          lpe0         = 1.8e-007          
+llpe0        = 1.1e-016          lpeb         = 0                 vbm          = -3                
+dvt0         = 1.14              ldvt0        = -6.124e-008       dvt1         = 0.22              
+ldvt1        = 2e-009            dvt2         = -0.02944          dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            dwg          = 0                 dwb          = 0
***************************************************************************                                                                                    
*             BASIC: Mobility Related Parameter                                                                                                                
***************************************************************************                                                                                    
+u0           = 0.028012+du0_n18_rf_mismatch                                                            
+lu0          = 5.4e-010+dlu0_n18_rf                                                           
+wu0          = -4.51e-010+dwu0_n18_rf                                                         
+pu0          = 4.6575e-016+dpu0_n18_rf                                                        
+ua           = -1.8869e-009      lua          = -3e-017           wua          = 7.6568e-017       
+pua          = 6.4915e-024       ub           = 3.515e-018        lub          = 2.92e-026         
+wub          = -1.274e-025       pub          = -7.86e-033        uc           = 1.4426e-010       
+luc          = 2.1688e-018       wuc          = -1.2768e-017      puc          = 8e-025            
+ud           = 0                 eu           = 1.67              
+vsat         = 70000+dvsat_n18_rf_mismatch                                                             
+lvsat        = 0.0006+dlvsat_n18_rf                                                           
+pvsat        = 5.2036e-010+dpvsat_n18_rf                                                      
+a0           = 1.6               la0          = -4e-007           pa0          = 5e-014            
+ags          = 0.56              lags         = 1.5e-007          wags         = -3e-008           
+pags         = 6e-014            b0           = 0                 b1           = 0                 
+keta         = -0.045548         lketa        = -7.6454e-009      wketa        = 1.0136e-008       
+pketa        = -1e-015           a1           = 0                 a2           = 0.99                                                                         
***************************************************************************  
*             BASIC: Subthreshold Related Parameter                           
***************************************************************************    
+voff         = -0.15+dvoff_n18_rf                                                             
+pvoff        = -5e-016           voffl        = 0                 minv         = 0                 
+nfactor      = 1                 eta0         = 0.14              peta0        = -6e-016           
+etab         = -0.07             petab        = 3.6e-015          dsub         = 0.56              
+cit          = 0.00065           lcit         = 1.6e-010          pcit         = -1e-018           
+cdsc         = 0                 cdscb        = 0                 cdscd        = 0.0001
***************************************************************************                                                                                    
*             BASIC: Output Resistance Related Parameter                                                                                                       
***************************************************************************                                                                                    
+pclm         = 0.31747           ppclm        = 4e-015            pdiblc1      = 0.04              
+pdiblc2      = 0.002             pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 3.45e+008         pscbe2       = 1e-006            pvag         = 0                 
+delta        = 0.001             pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 lambda       = 0 
***************************************************************************                                                                                    
*             Asymmetric and Bias-Dependent                                                                                                                    
***************************************************************************                                                                                    
+rdsw         = 90                rdswmin      = 0                 rdw          = 47                
+rdwmin       = 0                 rsw          = 47                rswmin       = 0                 
+prwg         = 0                 prwb         = 0                 wr           = 1  
***************************************************************************                                                                                    
*             Impact Ionization Current Model Parameters                                                                                                       
***************************************************************************                                                                                    
+alpha0       = 0                 alpha1       = 4.1739            lalpha1      = 2e-007            
+walpha1      = 4.64e-008         palpha1      = 2.5e-014          beta0        = 15.901    
***************************************************************************                                                                                    
*             Gate Dielectric Tunneling Current                                                                                                                
***************************************************************************                                                                                    
+aigbacc      = 0.43              bigbacc      = 0.054             cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0088021         bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.015123          bigc         = 0.0017647         cigc         = 0.0702            
+dlcig        = 1e-012            aigsd        = 0.0038304         waigsd       = -2e-010           
+paigsd       = -5e-018           bigsd        = 0.00030435        cigsd        = 0.19301           
+nigc         = 1.288             poxedge      = 1                 pigcd        = 1                 
+ntox         = 1                 toxref       = 3e-009          
***************************************************************************                                                                                    
*             GIDL Effect Parameters                                                                                                                           
***************************************************************************                                                                                    
+agidl        = 8.5074e-007       wagidl       = 2e-013            bgidl        = 2.9037e+009       
+wbgidl       = -50               cgidl        = 0.1               egidl        = 0.1        
***************************************************************************                                                                                    
*             Flicker Noise Model Parameter                                                                                                                    
***************************************************************************                                                                                    
+noia         = 6.24173e+041      noib         = 1.42569e+022      noic         = 6.62e+008                                                                    
+em           = 54761.2           ef           = 0.98              lintnoi      = -2e-008                                                                      
+ntnoi        = 1 
***************************************************************************                                                                                    
*             High-Speed RF Model Parameters                                                                                                                   
***************************************************************************                                                                                    
+rnoia=(-2.6579E-01*log(lrr)-3.3425E+00) tnoia=(1.8380E+06*log(lrr)+3.1801E+07) rnoib=0 tnoib=2e6                                                                                                                                                                
***************************************************************************                                                                                    
*             Capacitance Parameter                                                                                                                            
***************************************************************************                                                                                    
+xpart        = 0                                                                                                                                              
+cgdo         = 1.8e-010+dcgdo_n18_rf                                                                                                                        
+cgso         = 1.8e-010+dcgdo_n18_rf                                                                                                                        
+cgbo         = 0                                                                                                                                              
+cgdl         = 9e-011*kcgdl+dcgdl_n18_rf                                                                                                                          
+cgsl         = 9e-011*kcgdl+dcgdl_n18_rf                                                                                                                          
+cf           = (8.54e-011+dcf_n18_rf)                                                                                                                         
+clc          = 0                 cle          = 0.6               dlc          = 2.8339e-008*kdlc                                                                  
+dwc          = 0                 vfbcv        = -1                noff         = 1.6804                                                                       
+lnoff        = 1e-007            voffcv       = -0.020304         lvoffcv      = -2.088e-009                                                                  
+acde         = 0.384             moin         = 8                                                                                                       

*+dwc          = 0                 vfbcv        = -1                noff         = 1.6804                                                                     
*+lnoff        = 1e-007            voffcv       = -0.015        lvoffcv      = 0   
*+lnoff        = 1e-007            voffcv       = -0.02        lvoffcv      = 0                                                                
                                                             
*************************************************************************** 
*             Souce|Drain Junction Diode Model Parameter                     
***************************************************************************   
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.5              jss          = 1.1508e-006       jsws         = 1.4205e-014       
+jswgs        = 1.134e-013        jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 2e-008            
+jtsswgd      = 6e-009            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                                                                                                                                               
+cjs          = 0                                                                                                                        
+cjsws        = 0                                                                                                                     
+cjswgs       = 0                                                                                                                    
+mjs          = 0.34744           mjsws        = 0.19672           mjswgs       = 0.84898           
+pbs          = 0.70413           pbsws        = 0.58719           pbswgs       = 1.6255                                                                                                                                                               
***************************************************************************                                                                                    
*             Temperature coefficient                                                                                                                          
***************************************************************************                                                                                    
+tnom         = 25                ute          = -1.4012           lute         = 1.48e-008         
+kt1          = -0.24949          kt1l         = -2.9274e-009      kt2          = -0.05             
+wkt2         = 4e-009            ua1          = 1.76e-009         wua1         = -1.1e-016         
+pua1         = 1.625e-023        ub1          = -1.9392e-018      lub1         = -8.232e-026       
+wub1         = 1e-026            pub1         = -3.12e-033        uc1          = 1.124e-010        
+luc1         = -1.62e-017        puc1         = -3e-024           at           = 31820             
+pat          = -2.1e-010         prt          = 0                 njs          = 1.1294            
+xtis         = 3                 tpb          = 0.001             tpbsw        = 0.000868          
+tpbswg       = 0.0015811         tcj          = 0.00083836        tcjsw        = 0.0014935         
+tcjswg       = 0.0006583         tvoff        = 0                                                                                                               
***************************************************************************                                                                                    
*             Stress Effect Related Parameter                                                                                                                  
***************************************************************************                                                                                    
+saref        = 4.48e-006         sbref        = 4.48e-006         wlod         = 0                 
+ku0          = -4.5e-008         kvsat        = 1                 tku0         = 0                 
+lku0         = 7e-007            wku0         = 5e-007            pku0         = 7e-013            
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 3.5e-009          
+lkvth0       = -6e-008           wkvth0       = 1e-007            pkvth0       = 2e-014            
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                                                                                                                                                                
***************************************************************************                                                                                    
*             Well Proximity Effect Model Parameters                                                                                                           
***************************************************************************                                                                                    
+web          = 0                 wec          = 0                 kvth0we      = 0                                                                            
+k2we         = 0                 ku0we        = 0                 scref        = 1e-006                                                                       
***rf***                                                                                                                                                       
+ XRCRG1  = 12              XRCRG2  = 1                                                                                                                      
+ RSHG    =(rshg_n18_rf)                                                                                                                                               
******************************************************
//* **
model ndio18_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 1.1508e-006 isw = 1.4205e-014 vb = 11.5 ibv = 55.6 
+n = 1.1294 ns = 1.1294 rs = 5.0328e-010 
+cj = 0.00098714+dcj_n18_rf cjsw = 5.8272e-011*0.7+dcjsw_n18_rf vj = 0.70413 vjsw = 0.58719 
+fcs = 0 mj = 0.34744 mjsw = 0.2 fc = 0 
+tlev = 1 tlevc = 1 trs = 0.0019296 xti = 3 
+cta = 0.00083836 ctp = 0.001 pta = 0.001395 ptp = 0.000868 
+eg = 1.16  tcv = -0.0004
* *                           
// **
model diobpw_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 1.0388e-006 isw = 1.4035e-013 vb = 15.5 ibv = 55.6 
+n = 1.1225 ns = 1.1225 rs = 1.8727e-010 
+cj = 0.00049858+dcj_diobpw_rf cjsw = 3.9867e-010+dcjsw_diobpw_rf vj = 0.67589 vjsw = 0.88873 
+fcs = 0 mj = 0.33041 mjsw = 0.444 fc = 0 
+tlev = 1 tlevc = 1 trs = 0.00035608 xti = 3 
+cta = 0.00090633 ctp = 0.00080455 pta = 0.001448 ptp = 0.0012196 
+eg = 1.16  tcv = -0.0005
// **
model dnwdio_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 2.1632e-006 isw = 1.177e-012 vb = 16 ibv = 55.556 
+n = 1.0435 ns = 1.0435 rs = 1.3973e-007 
+cj = 0.00013824+dcj_dnwdio_rf cjsw = 4.1094e-010+dcjsw_dnwdio_rf vj = 0.52465 vjsw = 0.62598 
+fcs = 0 mj = 0.32294 mjsw = 0.35115 fc = 0 
+tlev = 1 tlevc = 1 trs = 1e-005 xti = 3 
+cta = 0.001326 ctp = 0.001221 pta = 0.0013127 ptp = 0.0015078 
+eg = 1.16 gap1 = 7.02e-04 tcv = -0.0006
// *

ends dnw18_6t_ckt_rf_r


// *1.8v pmos (tt corner)
// * 1=drain,2=gate,3=source,4=bulk
inline subckt p18_ckt_rf_r (1 2 3 4)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 
//*****************************************
+Cgd_rf = (((0.4477e-15*(wrr*1e+6)**0.7545+0.1652e-15)*(lrr*1e+6)**0.36+(-0.3216e-15*(wrr*1e+6)**0.6796+0.2989e-15))*nfr)
+Cgs_rf = (((0.144e-15*(wrr*1e+6)**0.6414+0.3587e-15)*(lrr*1e+6)**0.36+(-0.171e-15*(wrr*1e+6)**0.664+0.2733e-15))*nfr+1.2e-15)
+Rg_rf = (((91.5*(wrr*1e+6)**-1.6+1.2)*(lrr*1e+6)**-1)*(nfr+6)**-1*0.75)
+Rsub1_rf = (200/nfr)
+Rsub2_rf = (((268.7*(wrr*1e+6)**-0.5+77.85)*(lrr*1e+6)**-1-286.8)*(nfr+4)**-1)
+Djdb_AREA_rf = (int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6))
+Djdb_PJ_rf   = (int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*8.7477))
+Djsb_AREA_rf = (int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6)
+Djsb_PJ_rf   = (int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*8.7477))
//*****************************************
Lgate       (2 20)  inductor l=1e-12                        m=mrr
Rgate       (20 21) resistor r=(Rg_rf*(1+drg_p18_rf))       m=mrr
Cgd_ext     (21 11) capacitor c=(Cgd_rf*(1+dcgdext_p18_rf)) m=mrr
Cgs_ext     (21 31) capacitor c=(Cgs_rf*(1+dcgsext_p18_rf)) m=mrr
Cds_ext     (15 31) capacitor c=1e-18                       m=mrr
Rds         (11 15) resistor r=1e-3                         m=mrr
Ldrain       (1 11) inductor l=1e-12                        m=mrr
Lsource      (3 31) inductor l=1e-12                        m=mrr
//*****************************************
Djdb  (11 12) pdio18_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf     m=mrr
Djsb  (31 32) pdio18_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf     m=mrr
//*****************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
//*****************************************
p18_ckt_rf_r (11 21 31 41) p18_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model p18_ckt_r bsim4 type = p
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 1                 igbmod       = 1                 wpemod       = 0                 

***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 1.5e-007          lmax         = 0.0001            wmin         = 1.9e-007          
+wmax         = 0.0001
***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               
+toxe         = 4.27e-009+dtoxe_p18_mismatch_rf                                                
+dtox         = 4.49e-010         xj           = 1.6e-007          ndep         = 1.0196e+017       
+ngate        = 1.4e+020          nsd          = 1e+020            rsh          = 6.75              
***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 4e-015            wln          = 1                 ww           = -2.9e-015         
+wwn          = 1                 wwl          = -1.6e-021         ll           = 5.8e-015          
+lln          = 1                 lw           = -5e-015           lwn          = 1                 
+lwl          = 2.1e-022          llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 wint         = 8e-009            lint         = -3.8e-008  
***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                 
+xgw          = 0.31e-6                 xgl          = 0                 
+xl           = -1.3e-008+dxl_p18_rf                                                           
+xw           = 4.2e-008+dxw_p18_rf                                                            

***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = -0.424+dvth0_p18_mismatch_rf                                                             
+lvth0        = 6.0043e-009+dlvth0_p18_rf                                                       
+wvth0        = 7.0678e-009+dwvth0_p18_rf                                                       
+pvth0        = -2.5096e-015+dpvth0_p18_rf                                                      
+vfb          = -1                phin         = 0.00784           k1           = 0.59936           
+wk1          = -1.224e-008       pk1          = 4.864e-016        k2           = 0.001             
+lk2          = 1.6077e-009       k3           = 10                k3b          = -0.52             
+w0           = 9.0826e-006       
+lpe0         = 8.3442e-008+dlpe0_p18_rf                                                       
+llpe0        = -3.1e-015         lpeb         = 0                 vbm          = -3                
+dvt0         = 0.10912           dvt1         = 0.7               pdvt1        = -2e-014           
+dvt2         = -0.04             dvtp0        = 0                 dvtp1        = 0                 
+dvt0w        = 0                 dvt1w        = 5724000           dvt2w        = -0.032            
+dwg          = 0                 dwb          = 0   
***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.0095+du0_p18_mismatch_rf                                                     
+lu0          = 6.4546e-010+dlu0_p18_rf                                                           
+wu0          = -4.8639e-010+dwu0_p18_rf                                                       
+pu0          = -5.65e-017+dpu0_p18_rf                                                         
+ua           = 4.5895e-010       lua          = -5.1955e-017      wua          = -1.9101e-016      
+pua          = -8.5072e-024      ub           = 1.186e-018        lub          = 1.8e-025          
+wub          = -3.4e-026         pub          = -2.9e-032         uc           = -9e-013           
+luc          = 2.66e-017         wuc          = -3.1137e-017      puc          = -5e-024           
+ud           = 0                 eu           = 1                
+vsat         = 90000+dvsat_p18_mismatch_rf                                                    
+lvsat        = 0.017934+dlvsat_p18_rf                                                         
+pvsat        = -4.2733e-009+dpvsat_p18_rf                                                     
+a0           = 1.3               ags          = 0.36618           lags         = 1.5e-007          
+wags         = 2.4972e-008       pags         = -8e-014           b0           = 1.5e-008          
+b1           = 0                 keta         = -0.02492          lketa        = -1.3175e-009      
+wketa        = 2e-008            pketa        = -1.2e-015         a1           = 0                 
+a2           = 0.99  
***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.13138+dvoff_p18_mismatch_rf                                                 
+voffl        = 0                 
+minv         = 0+dminv_p18_rf                                                                 
+lminv        = 0+dlminv_p18_rf                                                                
+nfactor      = 1                 eta0         = 0.197             leta0        = -8e-009           
+peta0        = 1e-015            etab         = -0.16842          dsub         = 0.56              
+cit          = 0.0012            lcit         = 1.6e-010          pcit         = 4.5e-017          
+cdsc         = 0                 cdscb        = 0                 cdscd        = 0.0001 
***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.45942           pdiblc1      = 1e-006            pdiblc2      = 0.00316           
+lpdiblc2     = 1.4e-009          pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 3.45e+008         pscbe2       = 1e-006            pvag         = 0                 
+delta        = 0.0049056         pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 lambda       = 0 
***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 560               rdswmin      = 0                 rdw          = 0                 
+rdwmin       = 0                 rsw          = 280               rswmin       = 0                 
+prwg         = 0.4               prwb         = 0                 wr           = 1    
***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 1e-007            alpha1       = 6.3468            lalpha1      = 3.125e-007        
+walpha1      = 7.4012e-006       beta0        = 22.77             wbeta0       = 7.2864e-007    
***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.38872           bigbacc      = 0.056592          cigbacc      = 0.0726            
+nigbacc      = 1.112             aigbinv      = 0.0094803         bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.0092217         bigc         = 0.0019436         cigc         = 0.0702            
+dlcig        = 1e-012            aigsd        = 0.0029613         bigsd        = 0.00013888        
+cigsd        = 0.0786            nigc         = 1.288             poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 3e-009   
***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 1e-007            bgidl        = 2.7937e+009       pbgidl       = -2.2e-005         
+cgidl        = 0.2027            egidl        = 0.084       
***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 8e+041            noib         = 1.42569e+022      noic         = 1.20341e+010      
+em           = 54761.2           ef           = 1.1               lintnoi      = -3e-008           
+ntnoi        = 1 
***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_p18_rf)                     xrcrg1 = 10                       xrcrg2  = 3
+rnoia=(0.0485*log(lrr)+1.2694)     tnoia=116.6e6      rnoib=0        tnoib=2e6 
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 2.1e-010+dcgdo_p18_rf                                                          
+cgso         = 2.1e-010+dcgdo_p18_rf                                                          
+cgbo         = 0                 
+cgdl         = 1.761e-010+dcgdl_p18_rf                                                        
+cgsl         = 1.761e-010+dcgdl_p18_rf                                                        
+cf           = 8.5e-011+dcf_p18_rf                                                            
+clc          = 0                 cle          = 0.6               dlc          = 4.5009e-008       
+dwc          = 0                 vfbcv        = -1                noff         = 1.9376            
+lnoff        = 1.232e-007        voffcv       = -0.001            lvoffcv      = -6.728e-009       
+acde         = 0.57425           lacde        = -1.92e-008        moin         = 5                 

***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 10.8              jss          = 3.1581e-007       jsws         = 5.4158e-015       
+jswgs        = 1.7175e-013       jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 1e-011            
+jtsswgd      = 5e-009            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                  
+cjs          = 0                                                           
+cjsws        = 0                                                       
+cjswgs       = 0                                                      
+mjs          = 0.41824           mjsws        = 0.2959            mjswgs       = 0.43777           
+pbs          = 0.79266           pbsws        = 0.76922           pbswgs       = 0.74096         
***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.049            lute         = -3e-008           
+wute         = 3e-008            kt1          = -0.27376          kt1l         = -8.3e-009         
+kt2          = -0.04384          ua1          = 1.76e-009         lua1         = -7.62e-017        
+wua1         = -8.0657e-017      pua1         = -5.64e-025        ub1          = -3.2196e-018      
+lub1         = -1.6264e-025      wub1         = 3.1968e-025       pub1         = 3.6e-032          
+uc1          = -1e-010           luc1         = 5.848e-018        wuc1         = 3e-017            
+puc1         = -3.5839e-024      at           = 500               pat          = -1.776e-009       
+prt          = 0                 njs          = 1.0918            xtis         = 3                 
+tpb          = 0.00038165        tpbsw        = 0.0009004         tpbswg       = 0.0020341         
+tcj          = 0.00084383        tcjsw        = 0.0014196         tcjswg       = 0.00088262        
+tvoff        = 0   
***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 4.48e-006         sbref        = 4.48e-006         wlod         = 0                 
+ku0          = 8e-008            kvsat        = -1                tku0         = 0                 
+lku0         = 1.5e-007          wku0         = 0                 pku0         = 2e-014            
+llodku0      = 1                 wlodku0      = 1                 kvth0        = -1e-010           
+lkvth0       = -1e-007           wkvth0       = -2e-007           pkvth0       = 2e-014            
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1
***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 0                 wec          = 0                 kvth0we      = 0                 
+k2we         = 0                 ku0we        = 0                 scref        = 1e-006            
*****************************************************************************   
// *
model pdio18_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 4e-010 perim = 8e-005 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 9.5099e-008 isw = 2.9999e-014 vb = 10.6 ibv = 2500 
+n = 0.99836 ns = 0.99836 rs = 3.6817e-010 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = (0.001*(1+dcj_pdio18_rf)) cjp = (8.0e-011*(1+dcjp_pdio18_rf)) vj = 0.84022 vjsw = 0.43076 
+fcs = 0 mj = 0.31824 mjsw = 0.21959 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 trs = 0.0022422 xti = 3 
+cta = 0.0010193 ctp = 0.00040931 pta = 0.0014196 ptp = 0.0009004 
+eg = 1.16 


ends p18_ckt_rf




// *1.8v pmos with psub as 5th terminal
// * 1=drain,2=gate,3=source,4=bulk,5=psub
inline subckt p18_5t_ckt_rf_r (1 2 3 4 5)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 arnwr=1e-12 pjnwr=4e-6
//*****************************************
+Cgd_rf = (((0.4477e-15*(wrr*1e+6)**0.7545+0.1652e-15)*(lrr*1e+6)**0.36+(-0.3216e-15*(wrr*1e+6)**0.6796+0.2989e-15))*nfr)
+Cgs_rf = (((0.144e-15*(wrr*1e+6)**0.6414+0.3587e-15)*(lrr*1e+6)**0.36+(-0.171e-15*(wrr*1e+6)**0.664+0.2733e-15))*nfr+1.2e-15)
+Rg_rf = (((91.5*(wrr*1e+6)**-1.6+1.2)*(lrr*1e+6)**-1)*(nfr+6)**-1*0.75)
+Rsub1_rf = (200/nfr)
+Rsub2_rf = (((268.7*(wrr*1e+6)**-0.5+77.85)*(lrr*1e+6)**-1-286.8)*(nfr+4)**-1)
+Djdb_AREA_rf = (int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6))
+Djdb_PJ_rf   = (int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*8.7477))
+Djsb_AREA_rf = (int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6)
+Djsb_PJ_rf   = (int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*8.7477))
//*****************************************
Lgate       (2 20)  inductor l=1e-12                        m=mrr
Rgate       (20 21) resistor r=(Rg_rf*(1+drg_p18_rf))       m=mrr
Cgd_ext     (21 11) capacitor c=(Cgd_rf*(1+dcgdext_p18_rf)) m=mrr
Cgs_ext     (21 31) capacitor c=(Cgs_rf*(1+dcgsext_p18_rf)) m=mrr
Cds_ext     (15 31) capacitor c=1e-18                       m=mrr
Rds         (11 15) resistor r=1e-3                         m=mrr
Ldrain       (1 11) inductor l=1e-12                        m=mrr
Lsource      (3 31) inductor l=1e-12                        m=mrr
//*****************************************
Djdb  (11 12) pdio18_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf     m=mrr
Djsb  (31 32) pdio18_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf     m=mrr
Djnw  (5 4)   nwdio_rf  AREA=arnwr PJ=pjnwr                 m=mrr 
//*****************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
//*****************************************
p18_5t_ckt_rf_r (11 21 31 41) p18_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model p18_ckt_r bsim4 type = p
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 1                 igbmod       = 1                 wpemod       = 0                 

***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 1.5e-007          lmax         = 0.0001            wmin         = 1.9e-007          
+wmax         = 0.0001
***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               
+toxe         = 4.27e-009+dtoxe_p18_mismatch_rf                                                
+dtox         = 4.49e-010         xj           = 1.6e-007          ndep         = 1.0196e+017       
+ngate        = 1.4e+020          nsd          = 1e+020            rsh          = 6.75              
***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 4e-015            wln          = 1                 ww           = -2.9e-015         
+wwn          = 1                 wwl          = -1.6e-021         ll           = 5.8e-015          
+lln          = 1                 lw           = -5e-015           lwn          = 1                 
+lwl          = 2.1e-022          llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 wint         = 8e-009            lint         = -3.8e-008  
***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                 
+xgw          = 0.31e-6                 xgl          = 0                 
+xl           = -1.3e-008+dxl_p18_rf                                                           
+xw           = 4.2e-008+dxw_p18_rf                                                            

***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = -0.424+dvth0_p18_mismatch_rf                                                             
+lvth0        = 6.0043e-009+dlvth0_p18_rf                                                       
+wvth0        = 7.0678e-009+dwvth0_p18_rf                                                       
+pvth0        = -2.5096e-015+dpvth0_p18_rf                                                      
+vfb          = -1                phin         = 0.00784           k1           = 0.59936           
+wk1          = -1.224e-008       pk1          = 4.864e-016        k2           = 0.001             
+lk2          = 1.6077e-009       k3           = 10                k3b          = -0.52             
+w0           = 9.0826e-006       
+lpe0         = 8.3442e-008+dlpe0_p18_rf                                                       
+llpe0        = -3.1e-015         lpeb         = 0                 vbm          = -3                
+dvt0         = 0.10912           dvt1         = 0.7               pdvt1        = -2e-014           
+dvt2         = -0.04             dvtp0        = 0                 dvtp1        = 0                 
+dvt0w        = 0                 dvt1w        = 5724000           dvt2w        = -0.032            
+dwg          = 0                 dwb          = 0   
***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.0095+du0_p18_mismatch_rf                                                     
+lu0          = 6.4546e-010+dlu0_p18_rf                                                           
+wu0          = -4.8639e-010+dwu0_p18_rf                                                       
+pu0          = -5.65e-017+dpu0_p18_rf                                                         
+ua           = 4.5895e-010       lua          = -5.1955e-017      wua          = -1.9101e-016      
+pua          = -8.5072e-024      ub           = 1.186e-018        lub          = 1.8e-025          
+wub          = -3.4e-026         pub          = -2.9e-032         uc           = -9e-013           
+luc          = 2.66e-017         wuc          = -3.1137e-017      puc          = -5e-024           
+ud           = 0                 eu           = 1                
+vsat         = 90000+dvsat_p18_mismatch_rf                                                    
+lvsat        = 0.017934+dlvsat_p18_rf                                                         
+pvsat        = -4.2733e-009+dpvsat_p18_rf                                                     
+a0           = 1.3               ags          = 0.36618           lags         = 1.5e-007          
+wags         = 2.4972e-008       pags         = -8e-014           b0           = 1.5e-008          
+b1           = 0                 keta         = -0.02492          lketa        = -1.3175e-009      
+wketa        = 2e-008            pketa        = -1.2e-015         a1           = 0                 
+a2           = 0.99  
***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.13138+dvoff_p18_mismatch_rf                                                 
+voffl        = 0                 
+minv         = 0+dminv_p18_rf                                                                 
+lminv        = 0+dlminv_p18_rf                                                                
+nfactor      = 1                 eta0         = 0.197             leta0        = -8e-009           
+peta0        = 1e-015            etab         = -0.16842          dsub         = 0.56              
+cit          = 0.0012            lcit         = 1.6e-010          pcit         = 4.5e-017          
+cdsc         = 0                 cdscb        = 0                 cdscd        = 0.0001 
***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.45942           pdiblc1      = 1e-006            pdiblc2      = 0.00316           
+lpdiblc2     = 1.4e-009          pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 3.45e+008         pscbe2       = 1e-006            pvag         = 0                 
+delta        = 0.0049056         pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 lambda       = 0 
***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 560               rdswmin      = 0                 rdw          = 0                 
+rdwmin       = 0                 rsw          = 280               rswmin       = 0                 
+prwg         = 0.4               prwb         = 0                 wr           = 1    
***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 1e-007            alpha1       = 6.3468            lalpha1      = 3.125e-007        
+walpha1      = 7.4012e-006       beta0        = 22.77             wbeta0       = 7.2864e-007    
***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.38872           bigbacc      = 0.056592          cigbacc      = 0.0726            
+nigbacc      = 1.112             aigbinv      = 0.0094803         bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.0092217         bigc         = 0.0019436         cigc         = 0.0702            
+dlcig        = 1e-012            aigsd        = 0.0029613         bigsd        = 0.00013888        
+cigsd        = 0.0786            nigc         = 1.288             poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 3e-009   
***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 1e-007            bgidl        = 2.7937e+009       pbgidl       = -2.2e-005         
+cgidl        = 0.2027            egidl        = 0.084       
***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 8e+041            noib         = 1.42569e+022      noic         = 1.20341e+010      
+em           = 54761.2           ef           = 1.1               lintnoi      = -3e-008           
+ntnoi        = 1 
***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_p18_rf)                     xrcrg1 = 10                       xrcrg2  = 3
+rnoia=(0.0485*log(lrr)+1.2694)     tnoia=116.6e6      rnoib=0        tnoib=2e6 
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 2.1e-010+dcgdo_p18_rf                                                          
+cgso         = 2.1e-010+dcgdo_p18_rf                                                          
+cgbo         = 0                 
+cgdl         = 1.761e-010+dcgdl_p18_rf                                                        
+cgsl         = 1.761e-010+dcgdl_p18_rf                                                        
+cf           = 8.5e-011+dcf_p18_rf                                                            
+clc          = 0                 cle          = 0.6               dlc          = 4.5009e-008       
+dwc          = 0                 vfbcv        = -1                noff         = 1.9376            
+lnoff        = 1.232e-007        voffcv       = -0.001            lvoffcv      = -6.728e-009       
+acde         = 0.57425           lacde        = -1.92e-008        moin         = 5                 

***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 10.8              jss          = 3.1581e-007       jsws         = 5.4158e-015       
+jswgs        = 1.7175e-013       jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 1e-011            
+jtsswgd      = 5e-009            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                  
+cjs          = 0                                                           
+cjsws        = 0                                                       
+cjswgs       = 0                                                      
+mjs          = 0.41824           mjsws        = 0.2959            mjswgs       = 0.43777           
+pbs          = 0.79266           pbsws        = 0.76922           pbswgs       = 0.74096         
***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.049            lute         = -3e-008           
+wute         = 3e-008            kt1          = -0.27376          kt1l         = -8.3e-009         
+kt2          = -0.04384          ua1          = 1.76e-009         lua1         = -7.62e-017        
+wua1         = -8.0657e-017      pua1         = -5.64e-025        ub1          = -3.2196e-018      
+lub1         = -1.6264e-025      wub1         = 3.1968e-025       pub1         = 3.6e-032          
+uc1          = -1e-010           luc1         = 5.848e-018        wuc1         = 3e-017            
+puc1         = -3.5839e-024      at           = 500               pat          = -1.776e-009       
+prt          = 0                 njs          = 1.0918            xtis         = 3                 
+tpb          = 0.00038165        tpbsw        = 0.0009004         tpbswg       = 0.0020341         
+tcj          = 0.00084383        tcjsw        = 0.0014196         tcjswg       = 0.00088262        
+tvoff        = 0   
***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 4.48e-006         sbref        = 4.48e-006         wlod         = 0                 
+ku0          = 8e-008            kvsat        = -1                tku0         = 0                 
+lku0         = 1.5e-007          wku0         = 0                 pku0         = 2e-014            
+llodku0      = 1                 wlodku0      = 1                 kvth0        = -1e-010           
+lkvth0       = -1e-007           wkvth0       = -2e-007           pkvth0       = 2e-014            
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1
***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 0                 wec          = 0                 kvth0we      = 0                 
+k2we         = 0                 ku0we        = 0                 scref        = 1e-006            
*****************************************************************************      
// *
model pdio18_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 4e-010 perim = 8e-005 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 9.5099e-008 isw = 2.9999e-014 vb = 10.6 ibv = 2500 
+n = 0.99836 ns = 0.99836 rs = 3.6817e-010 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = (0.001*(1+dcj_pdio18_rf)) cjp = (8.0e-011*(1+dcjp_pdio18_rf)) vj = 0.84022 vjsw = 0.43076 
+fcs = 0 mj = 0.31824 mjsw = 0.21959 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 trs = 0.0022422 xti = 3 
+cta = 0.0010193 ctp = 0.00040931 pta = 0.0014196 ptp = 0.0009004 
+eg = 1.16 
//
model nwdio_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 9.6e-009 perim = 4e-004 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 2.3733e-006 isw = 2.9142e-014 vb = 15 ibv = 104 
+n = 1.085 ns = 1.085 rs = 8.4602e-009 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = (0.000131*(1+dcj_nwdio_rf)) cjp = (5.0047e-010*(1+dcjp_nwdio_rf)) vj = 0.41624 vjsw = 0.81575 
+fcs = 0 mj = 0.26295 mjsw = 0.377 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 trs = 0.0004 xti = 3 
+cta = 0.0017608 ctp = 0.0012659 pta = 0.00155 ptp = 0.0022128 
+eg = 1.16 
// *


ends p18_5t_ckt_rf


* 3.3v nmos 
* 1=drain,2=gate,3=source,4=bulk
inline subckt n33_ckt_rf_r (1 2 3 4)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 
**********************************************
+Rg_rf	       = max((1/(1.472E-32*pwr(lrr,-4.885)+0.497))*((1.987*exp(-5.279E+06*lrr))*(((0.0007874+51.24*wrr)+((-97.72)+(-5.316E7)*wrr)*lrr)+((5.049E-6+1.042*wrr)+((-3.595)+1.26E5*wrr)*lrr)*nfr)/wrr/nfr),1e-3)
+Cgd_rf        = max((1/(4.343e-11*pwr(lrr,-1.473)+0.97))*((0.0001332*lrr-2.01E-11)*wrr+(5.532E-12*lrr+4.606E-16))*nfr,1e-18)
+Cgs_rf	       = max((4.383E-43*pwr(lrr,-6.406)+0.99988)*(1.008*exp(-416800*wrr)+0.084)*(3.936e-16*log(lrr)+6.428E-15)*EXP(wrr*(-3.91224E11*lrr+195609))*nfr,1e-18)
+Cds_rf	       = 0.5*max((1.405e-11*pwr(wrr,-1.732)+0.797)*((-8.212e-11*log(lrr)-1.005e-9)*wrr-(1/(7.619E-18*pwr(lrr,-2.45)+0.179)*1e-17))*nfr,1e-18)

+Rsub1_rf      = max(-1.076E+08*lrr+256,1e-3)
+Rsub2_rf      = 0.01*max((((2.191E4+(-2.115E9)*wrr))+(((-428.3)+4.045E7*wrr))*nfr)/nfr,1e-3)
+Rsub3_rf      =  Rsub2_rf
+Rdc_n33_rf    = max((86.7923*exp(-0.1713*wrr*1e6)),1e-3)
+Rsc_n33_rf    = max((86.7923*exp(-0.1713*wrr*1e6)),1e-3)
+Rds_rf	       = max(460.31*exp(-223066*wrr),1e-3)
+Djdb_AREA_rf  = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf    = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)                                                                                          
+Djsb_AREA_rf  = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf    = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)  
**********************************************
Lgate       ( 2 20) inductor  l=1p                        m=mrr
Rgate       (20 21) resistor  r=Rg_rf*(1+drg_n33_rf)      m=mrr
Cgd_ext     (21 11) capacitor c=Cgd_rf*(1+dcgdext_n33_rf) m=mrr
Cgs_ext     (21 31) capacitor c=Cgs_rf*(1+dcgsext_n33_rf) m=mrr
Cds_ext     (15 31) capacitor c=Cds_rf                    m=mrr
Rds         (11 15) resistor  r=Rds_rf                    m=mrr
Ldrain       (1 11) inductor  l=1p                        m=mrr
Lsource      (3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (12 11) ndio33_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (32 31) ndio33_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
**********************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
**********************************************
n33_ckt_rf_r (11 21 31 41) n33_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model n33_ckt_r bsim4 type = n
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 0                 igbmod       = 0                 wpemod       = 0                 

***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 3.5e-007          lmax         = 0.0001            wmin         = 2.2e-007          
+wmax         = 0.0001            

***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               toxe         = 6.65e-009+dtoxe_n33_mismatch_rf         
+dtox         = 3.9e-010                                                          
+xj           = 1.6e-007          ndep         = 6.250661e+017     ngate        = 1.6e+020          
+rsh          = 12                

***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 1.02e-014         wln          = 1                 ww           = -2.677213e-015    
+wwn          = 1                 wwl          = -2.5e-021         ll           = -9.5e-015         
+lln          = 1                 lw           = 0                 lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 

***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                 
+xgw          = 0.31e-006                 xgl          = -1.38e-008                 
+xl           = -1.38e-008+dxl_n33_mismatch_rf                                                          
+xw           = 1.58e-008+dxw_n33_mismatch_rf                                                           

***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = 0.75619+dvth0_n33_mismatch_rf                                                           
+lvth0        = 2.0644e-009+dlvth0_n33_rf                                                      
+wvth0        = -1.6313e-008+dwvth0_n33_rf                                                     
+pvth0        = 2.393452e-015+dpvth0_n33_rf                                                    
+phin         = 0.15              k1           = 0.92              k2           = 0.0192267         
+lk2          = -1.7175e-008      wk2          = 1e-009            pk2          = 1.2125e-015       
+k3           = -1                lk3          = 3.247781e-006     wk3          = 1.174813e-006     
+pk3          = -2.895674e-013    k3b          = 2.7               lk3b         = -4.94e-006        
+wk3b         = 1.02e-006         pk3b         = 8.05e-013         w0           = 1.25e-006         
+lpe0         = 1.793508e-007     llpe0        = -3e-014           wlpe0        = -1.83375e-014     
+plpe0        = 2.8e-021          lpeb         = 0                 llpeb        = -1e-014           
+vbm          = -3                dvt0         = 1.977453          dvt1         = 0.81669           
+wdvt1        = 4.9e-009          dvt2         = -1.52658          dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            wint         = 3.409374e-008     lint         = 8.591858e-008     
+dwg          = -1e-009           wdwg         = 2.5e-016          dwb          = 0                 

***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.034389+du0_n33_mismatch_rf                                                            
+lu0          = -6.5037e-010+dlu0_n33_rf                                                       
+wu0          = 2.9719e-010+dwu0_n33_rf                                                        
+pu0          = 1.3e-016+dpu0_n33_rf                                                           
+ua           = -1.319673e-009    lua          = -3e-017           wua          = 4.255033e-017     
+pua          = -1.2e-023         ub           = 3.076021e-018     wub          = -1.578187e-025    
+pub          = 2e-033            uc           = 1.75496e-010      luc          = -6e-018           
+wuc          = -2e-017           puc          = -6e-025           ud           = 0                 
+eu           = 1.67              
+vsat         = 54975.69+dvsat_n33_mismatch_rf                                                          
+lvsat        = 0.0050622+dlvsat_n33_rf                                                        
+wvsat        = 0.001842913+dwvsat_n33_rf                                                      
+pvsat        = 1.370232e-010+dpvsat_n33_rf                                                    
+a0           = 1.446797          la0          = -3.3e-007         pa0          = 7e-014            
+ags          = 0.289501          lags         = 2.9e-007          wags         = -1.251297e-008    
+pags         = -1e-014           b0           = 8.604318e-008     lb0          = -6.913192e-014    
+wb0          = -4.812935e-014    pb0          = -1.044909e-020    b1           = 0                 
+lb1          = -1.606808e-014    wb1          = 1.713014e-013     pb1          = 8.347455e-021     
+keta         = -0.030075         lketa        = 1.391934e-009     pketa        = -7.784875e-015    
+a1           = 0                 a2           = 1                 

***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.147398+dvoff_n33_mismatch_rf         
+voffl        = -4.2e-009         minv         = -0.45             
+nfactor      = 1.066459          pnfactor     = -7e-015           eta0         = 0.08              
+etab         = -0.07             letab        = -1.7e-007         petab        = 2.5e-014          
+dsub         = 0.56              cit          = 4.634146e-005     cdsc         = 0.00024           
+cdscb        = 0                 cdscd        = 2e-005            

***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.26              pdiblc1      = 0.39              pdiblc2      = 0.000705          
+ppdiblc2     = -2.5e-017         pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 4.24e+008         pscbe2       = 1e-005            pvag         = 0                 
+delta        = 0                 ldelta       = 2e-009            fprout       = 0                 
+pdits        = 0                 pditsl       = 0                 pditsd       = 0                 

***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 549.89337         rdw          = 24                rdwmin       = 0                 
+rsw          = 24                rswmin       = 0                 prwg         = 0.108             
+prwb         = 0                 wr           = 1                 

***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 0                 alpha1       = 11.09775          lalpha1      = 2.123369e-005     
+beta0        = 25.056188         lbeta0       = 2e-006            

***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.002249          bigbacc      = 1.71e-007         cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0111            bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.00525           laigc        = -1.3e-010         waigc        = -1.2e-010         
+bigc         = 0.0003            cigc         = 0.075             dlcig        = 4e-009            
+aigsd        = 0.0045            waigsd       = -1e-010           bigsd        = 0.0001            
+cigsd        = 0.075             nigc         = 1                 poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 6.65e-009         

***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 0                 
+lagidl       = 0+dlagidl_n33_rf                                                               
+pagidl       = 0+dpagidl_n33_rf                                                               
+bgidl        = 2.3e+009          cgidl        = 0.5               egidl        = 0.8               

***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 6.25e+041         noib         = 5E+25        noic         = 8.75              
+em           = 4.1e+007          ef           = 1                 lintnoi      = 0                 
+ntnoi        = 1                 

***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_n33_rf)                     xrcrg1 = 10                       xrcrg2  = 8
+ngcon= 2
+rnoia = (max(0.01303+6.337*pwr(exp(10*(lrr*1e+6)),-0.8695)+0.56*pwr((wrr*1e+6),0.138),0.1))    tnoia = 0.1e+7    rnoib=0    tnoib=1.0e+7
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 1e-010+dcgdo_n33_rf                                                            
+cgso         = 1e-010+dcgso_n33_rf                                                            
+cgbo         = 0                 
+cgdl         = (2.6e-010+dcgdl_n33_rf)*0.8                                                          
+cgsl         = (2.6e-010+dcgsl_n33_rf)*0.8                                                          
+cf           = 7.55e-011+dcf_n33_rf
+clc          = 1e-007            cle          = 0.6               dlc          = 5.381e-008*(0.123*EXP(1404000*lr)+1)       
+dwc          = 0                 noff         = 2.2               lnoff        = 3.856e-007        
+voffcv       = -0.1184           lvoffcv      = -2.968e-008       acde         = 0.23814           
+moin         = 5.2               

***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.8              jss          = 4.1904e-007       jsws         = 3.9508e-013       
+jswgs        = 4.3285e-014       jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 
+jtsswgs      = 1.61e-009+djtsswgs_n33_rf                                                      
+jtsswgd      = 1.61e-009+djtsswgd_n33_rf                                                      
+njts         = 20                njtssw       = 20                njtsswg      = 20                
+xtss         = 0.02              xtsd         = 0.02              xtssws       = 0.02              
+xtsswd       = 0.02              xtsswgs      = 0.02              xtsswgd      = 0.02              
+vtss         = 10                vtsd         = 10                vtssws       = 10                
+vtsswd       = 10                vtsswgs      = 10                vtsswgd      = 10                
+tnjts        = 0               tnjtssw      = 0                 tnjtsswg     = 0                 
+cjs          = 0                                                        
+cjsws        = 0                                                      
+cjswgs       = 0                                                    
+mjs          = 0.32174           mjsws        = 0.0001727         mjswgs       = 0.36511           
+pbs          = 0.70384           pbsws        = 0.44462           pbswgs       = 0.59056           

***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.5              kt1          = -0.2565           
+lkt1         = 6e-009            pkt1         = 1.5e-015          kt2          = -0.0572           
+ua1          = 1e-009            ub1          = -1.29e-018        lub1         = -1e-025           
+wub1         = -1.17e-025        pub1         = 5e-032            uc1          = 5.6e-011          
+wuc1         = -1.68e-017        at           = 100000            lat          = -0.0157           
+pat          = 3e-010            njs          = 1.0296            xtis         = 3                 
+tpb          = 0.0016752         tpbsw        = 0.0009385         tpbswg       = 0.001502          
+tcj          = 0.00093975        tcjsw        = 0.00046393        tcjswg       = 0.0011153         
+tvoff        = 0.002             

***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 5.33e-006         sbref        = 5.33e-006         wlod         = 0                 
+ku0          = -2e-008           kvsat        = 1                 tku0         = 0                 
+lku0         = 5e-007            wku0         = 1e-006            pku0         = 0                 
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 6e-009            
+lkvth0       = 2e-007            wkvth0       = -5e-008           pkvth0       = 0                 
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                 

***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 1                 wec          = 1                 kvth0we      = 0            
+k2we         = 0                 ku0we        = 0           scref        = 1e-006            
*****************************************************************************************
* **
model ndio33_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
+dcap = 2 area = 4e-10 perim = 0.00008 tnom = 25 
+js = 4.1904e-007  isw = 3.9508e-013  expli = 1e+020 
+n = 1.0296  ns = 1.0296 rs = 2.8395e-010 jtun = 0 jtunsw = 0 
+ntun = 30 ibv = 2.50e+03 vb = 11.8 
+cj = 0.00086098+dcj_ndio33_rf cjsw = (9.677e-011+dcjsw_ndio33_rf)*0.5 vj = 0.70384 vjsw = 0.44462 
+fcs = 0 mj = 0.32174 mjsw = 0.16049 fc = 0 
+tt = 0 
+tlev = 1 tlevc = 1 tcv = 0 trs = 0.00065303 
+xti = 3 xtitun = 3 cta = 0.00093975 ctp = 0.00046393 
+pta = 0.0016752 ptp = 0.0009385 eg = 1.16 gap1 = 0.000702 
+gap2 = 1108 ttt1 = 0 ttt2 = 0 tm1 = 0 
+tm2 = 0 

ends n33_ckt_rf_r


* 3.3v nmos in dnw with 4 ports
* 1=drain,2=gate,3=source,4=bulk
inline subckt dnw33_ckt_rf_r (1 2 3 4)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 
**********************************************
+Rg_rf	       = max((1/(1.472E-32*pwr(lrr,-4.885)+0.497))*((1.987*exp(-5.279E+06*lrr))*(((0.0007874+51.24*wrr)+((-97.72)+(-5.316E7)*wrr)*lrr)+((5.049E-6+1.042*wrr)+((-3.595)+1.26E5*wrr)*lrr)*nfr)/wrr/nfr),1e-3)
+Cgd_rf        = max((1/(4.343e-11*pwr(lrr,-1.473)+0.97))*((0.0001332*lrr-2.01E-11)*wrr+(5.532E-12*lrr+4.606E-16))*nfr,1e-18)
+Cgs_rf	       = max((4.383E-43*pwr(lrr,-6.406)+0.99988)*(1.008*exp(-416800*wrr)+0.084)*(3.936e-16*log(lrr)+6.428E-15)*EXP(wrr*(-3.91224E11*lrr+195609))*nfr,1e-18)
+Cds_rf	       = 0.5*max((1.405e-11*pwr(wrr,-1.732)+0.797)*((-8.212e-11*log(lrr)-1.005e-9)*wrr-(1/(7.619E-18*pwr(lrr,-2.45)+0.179)*1e-17))*nfr,1e-18)
+Rsub1_rf      = max(-1.076E+08*lrr+256,1e-3)
+Rsub2_rf      = 0.01*max((((2.191E4+(-2.115E9)*wrr))+(((-428.3)+4.045E7*wrr))*nfr)/nfr,1e-3)
+Rsub3_rf      =  Rsub2_rf
+Rdc_n33_rf    = max((86.7923*exp(-0.1713*wrr*1e6)),1e-3)
+Rsc_n33_rf    = max((86.7923*exp(-0.1713*wrr*1e6)),1e-3)
+Rds_rf	       = max(460.31*exp(-223066*wrr),1e-3)
+Djdb_AREA_rf  = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf    = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)                                                                                          
+Djsb_AREA_rf  = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf    = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)  
**********************************************
Lgate       ( 2 20) inductor  l=1p                        m=mrr
Rgate       (20 21) resistor  r=Rg_rf*(1+drg_n33_rf)      m=mrr
Cgd_ext     (21 11) capacitor c=Cgd_rf*(1+dcgdext_n33_rf) m=mrr
Cgs_ext     (21 31) capacitor c=Cgs_rf*(1+dcgsext_n33_rf) m=mrr
Cds_ext     (15 31) capacitor c=Cds_rf                    m=mrr
Rds         (11 15) resistor  r=Rds_rf                    m=mrr
Ldrain       (1 11) inductor  l=1p                        m=mrr
Lsource      (3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (12 11) ndio33_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (32 31) ndio33_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
**********************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
**********************************************
dnw33_ckt_rf_r (11 21 31 41) n33_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model n33_ckt_r bsim4 type = n
**********************************************************************************************                                                                            
*                              3.3V CORE NMOS MODEL                               *                                                                            
**********************************************************************************************                                                                            
* GENERAL PARAMETERS                                                                                                                                           
*                                                                                                                                                              
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 0                 igbmod       = 0                 wpemod       = 0                 

***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 3.5e-007          lmax         = 0.0001            wmin         = 2.2e-007          
+wmax         = 0.0001            

***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               toxe         = 6.65e-009+dtoxe_n33_mismatch_rf         
+dtox         = 3.9e-010                                                          
+xj           = 1.6e-007          ndep         = 6.250661e+017     ngate        = 1.6e+020          
+rsh          = 12                

***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 1.02e-014         wln          = 1                 ww           = -2.677213e-015    
+wwn          = 1                 wwl          = -2.5e-021         ll           = -9.5e-015         
+lln          = 1                 lw           = 0                 lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 

***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                 
+xgw          = 0.31e-006                 xgl          = -1.38e-008                 
+xl           = -1.38e-008+dxl_n33_mismatch_rf                                                          
+xw           = 1.58e-008+dxw_n33_mismatch_rf                                                           

***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = 0.75619+dvth0_n33_mismatch_rf                                                           
+lvth0        = 2.0644e-009+dlvth0_n33_rf                                                      
+wvth0        = -1.6313e-008+dwvth0_n33_rf                                                     
+pvth0        = 2.393452e-015+dpvth0_n33_rf                                                    
+phin         = 0.15              k1           = 0.92              k2           = 0.0192267         
+lk2          = -1.7175e-008      wk2          = 1e-009            pk2          = 1.2125e-015       
+k3           = -1                lk3          = 3.247781e-006     wk3          = 1.174813e-006     
+pk3          = -2.895674e-013    k3b          = 2.7               lk3b         = -4.94e-006        
+wk3b         = 1.02e-006         pk3b         = 8.05e-013         w0           = 1.25e-006         
+lpe0         = 1.793508e-007     llpe0        = -3e-014           wlpe0        = -1.83375e-014     
+plpe0        = 2.8e-021          lpeb         = 0                 llpeb        = -1e-014           
+vbm          = -3                dvt0         = 1.977453          dvt1         = 0.81669           
+wdvt1        = 4.9e-009          dvt2         = -1.52658          dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            wint         = 3.409374e-008     lint         = 8.591858e-008     
+dwg          = -1e-009           wdwg         = 2.5e-016          dwb          = 0                 

***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.034389+du0_n33_mismatch_rf                                                            
+lu0          = -6.5037e-010+dlu0_n33_rf                                                       
+wu0          = 2.9719e-010+dwu0_n33_rf                                                        
+pu0          = 1.3e-016+dpu0_n33_rf                                                           
+ua           = -1.319673e-009    lua          = -3e-017           wua          = 4.255033e-017     
+pua          = -1.2e-023         ub           = 3.076021e-018     wub          = -1.578187e-025    
+pub          = 2e-033            uc           = 1.75496e-010      luc          = -6e-018           
+wuc          = -2e-017           puc          = -6e-025           ud           = 0                 
+eu           = 1.67              
+vsat         = 54975.69+dvsat_n33_mismatch_rf                                                          
+lvsat        = 0.0050622+dlvsat_n33_rf                                                        
+wvsat        = 0.001842913+dwvsat_n33_rf                                                      
+pvsat        = 1.370232e-010+dpvsat_n33_rf                                                    
+a0           = 1.446797          la0          = -3.3e-007         pa0          = 7e-014            
+ags          = 0.289501          lags         = 2.9e-007          wags         = -1.251297e-008    
+pags         = -1e-014           b0           = 8.604318e-008     lb0          = -6.913192e-014    
+wb0          = -4.812935e-014    pb0          = -1.044909e-020    b1           = 0                 
+lb1          = -1.606808e-014    wb1          = 1.713014e-013     pb1          = 8.347455e-021     
+keta         = -0.030075         lketa        = 1.391934e-009     pketa        = -7.784875e-015    
+a1           = 0                 a2           = 1                 

***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.147398+dvoff_n33_mismatch_rf         
+voffl        = -4.2e-009         minv         = -0.45             
+nfactor      = 1.066459          pnfactor     = -7e-015           eta0         = 0.08              
+etab         = -0.07             letab        = -1.7e-007         petab        = 2.5e-014          
+dsub         = 0.56              cit          = 4.634146e-005     cdsc         = 0.00024           
+cdscb        = 0                 cdscd        = 2e-005            

***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.26              pdiblc1      = 0.39              pdiblc2      = 0.000705          
+ppdiblc2     = -2.5e-017         pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 4.24e+008         pscbe2       = 1e-005            pvag         = 0                 
+delta        = 0                 ldelta       = 2e-009            fprout       = 0                 
+pdits        = 0                 pditsl       = 0                 pditsd       = 0                 

***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 549.89337         rdw          = 24                rdwmin       = 0                 
+rsw          = 24                rswmin       = 0                 prwg         = 0.108             
+prwb         = 0                 wr           = 1                 

***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 0                 alpha1       = 11.09775          lalpha1      = 2.123369e-005     
+beta0        = 25.056188         lbeta0       = 2e-006            

***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.002249          bigbacc      = 1.71e-007         cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0111            bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.00525           laigc        = -1.3e-010         waigc        = -1.2e-010         
+bigc         = 0.0003            cigc         = 0.075             dlcig        = 4e-009            
+aigsd        = 0.0045            waigsd       = -1e-010           bigsd        = 0.0001            
+cigsd        = 0.075             nigc         = 1                 poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 6.65e-009         

***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 0                 
+lagidl       = 0+dlagidl_n33_rf                                                               
+pagidl       = 0+dpagidl_n33_rf                                                               
+bgidl        = 2.3e+009          cgidl        = 0.5               egidl        = 0.8               

***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 6.25e+041         noib         = 5E+25        noic         = 8.75              
+em           = 4.1e+007          ef           = 1                 lintnoi      = 0                 
+ntnoi        = 1                 

***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_n33_rf)                     xrcrg1 = 10                       xrcrg2  = 8
+ngcon= 2
+rnoia = (max(0.01303+6.337*pwr(exp(10*(lrr*1e+6)),-0.8695)+0.56*pwr((wrr*1e+6),0.138),0.1))    tnoia = 0.1e+7    rnoib=0    tnoib=1.0e+7
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 1e-010+dcgdo_n33_rf                                                            
+cgso         = 1e-010+dcgso_n33_rf                                                            
+cgbo         = 0                 
+cgdl         = (2.6e-010+dcgdl_n33_rf)*0.8                                                          
+cgsl         = (2.6e-010+dcgsl_n33_rf)*0.8                                                          
+cf           = 7.55e-011+dcf_n33_rf
+clc          = 1e-007            cle          = 0.6               dlc          = 5.381e-008*(0.123*EXP(1404000*lr)+1)       
+dwc          = 0                 noff         = 2.2               lnoff        = 3.856e-007        
+voffcv       = -0.1184           lvoffcv      = -2.968e-008       acde         = 0.23814           
+moin         = 5.2               

***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.8              jss          = 4.1904e-007       jsws         = 3.9508e-013       
+jswgs        = 4.3285e-014       jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 
+jtsswgs      = 1.61e-009+djtsswgs_n33_rf                                                      
+jtsswgd      = 1.61e-009+djtsswgd_n33_rf                                                      
+njts         = 20                njtssw       = 20                njtsswg      = 20                
+xtss         = 0.02              xtsd         = 0.02              xtssws       = 0.02              
+xtsswd       = 0.02              xtsswgs      = 0.02              xtsswgd      = 0.02              
+vtss         = 10                vtsd         = 10                vtssws       = 10                
+vtsswd       = 10                vtsswgs      = 10                vtsswgd      = 10                
+tnjts        = 0               tnjtssw      = 0                 tnjtsswg     = 0                 
+cjs          = 0                                                        
+cjsws        = 0                                                      
+cjswgs       = 0                                                    
+mjs          = 0.32174           mjsws        = 0.0001727         mjswgs       = 0.36511           
+pbs          = 0.70384           pbsws        = 0.44462           pbswgs       = 0.59056           

***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.5              kt1          = -0.2565           
+lkt1         = 6e-009            pkt1         = 1.5e-015          kt2          = -0.0572           
+ua1          = 1e-009            ub1          = -1.29e-018        lub1         = -1e-025           
+wub1         = -1.17e-025        pub1         = 5e-032            uc1          = 5.6e-011          
+wuc1         = -1.68e-017        at           = 100000            lat          = -0.0157           
+pat          = 3e-010            njs          = 1.0296            xtis         = 3                 
+tpb          = 0.0016752         tpbsw        = 0.0009385         tpbswg       = 0.001502          
+tcj          = 0.00093975        tcjsw        = 0.00046393        tcjswg       = 0.0011153         
+tvoff        = 0.002             

***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 5.33e-006         sbref        = 5.33e-006         wlod         = 0                 
+ku0          = -2e-008           kvsat        = 1                 tku0         = 0                 
+lku0         = 5e-007            wku0         = 1e-006            pku0         = 0                 
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 6e-009            
+lkvth0       = 2e-007            wkvth0       = -5e-008           pkvth0       = 0                 
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                 

***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 1                 wec          = 1                 kvth0we      = 0            
+k2we         = 0                 ku0we        = 0           scref        = 1e-006            
*****************************************************************************************
* **

model ndio33_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
+dcap = 2 area = 4e-10 perim = 0.00008 tnom = 25 
+js = 4.1904e-007  isw = 3.9508e-013  expli = 1e+020 
+n = 1.0296  ns = 1.0296 rs = 2.8395e-010 jtun = 0 jtunsw = 0 
+ntun = 30 ibv = 2.50e+03 vb = 11.8 
+cj = 0.00086098+dcj_ndio33_rf cjsw = (9.677e-011+dcjsw_ndio33_rf)*0.5 vj = 0.70384 vjsw = 0.44462 
+fcs = 0 mj = 0.32174 mjsw = 0.16049 fc = 0 
+tt = 0 
+tlev = 1 tlevc = 1 tcv = 0 trs = 0.00065303 
+xti = 3 xtitun = 3 cta = 0.00093975 ctp = 0.00046393 
+pta = 0.0016752 ptp = 0.0009385 eg = 1.16 gap1 = 0.000702 
+gap2 = 1108 ttt1 = 0 ttt2 = 0 tm1 = 0 
+tm2 = 0 

ends dnw33_ckt_rf_r


* 3.3v nmos in dnw with 6 ports
* 1=drain,2=gate,3=source,4=bulk,5=dnw,6=psub
inline subckt dnw33_6t_ckt_rf_r (1 2 3 4 5 6)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.04e-006 sbrr=1.04e-006 sdrr=0.54e-6 nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 arpwr=162.01e-12 pjpwr=55.12e-6 ardnwr=190.57e-12 pjdnwr=59.12e-6
**********************************************
+Rg_rf	       = max((1/(1.472E-32*pwr(lrr,-4.885)+0.497))*((1.987*exp(-5.279E+06*lrr))*(((0.0007874+51.24*wrr)+((-97.72)+(-5.316E7)*wrr)*lrr)+((5.049E-6+1.042*wrr)+((-3.595)+1.26E5*wrr)*lrr)*nfr)/wrr/nfr),1e-3)
+Cgd_rf        = max((1/(4.343e-11*pwr(lrr,-1.473)+0.97))*((0.0001332*lrr-2.01E-11)*wrr+(5.532E-12*lrr+4.606E-16))*nfr,1e-18)
+Cgs_rf	       = max((4.383E-43*pwr(lrr,-6.406)+0.99988)*(1.008*exp(-416800*wrr)+0.084)*(3.936e-16*log(lrr)+6.428E-15)*EXP(wrr*(-3.91224E11*lrr+195609))*nfr,1e-18)
+Cds_rf	       = 0.5*max((1.405e-11*pwr(wrr,-1.732)+0.797)*((-8.212e-11*log(lrr)-1.005e-9)*wrr-(1/(7.619E-18*pwr(lrr,-2.45)+0.179)*1e-17))*nfr,1e-18)
+Rsub1_rf      = max(-1.076E+08*lrr+256,1e-3)
+Rsub2_rf      = 0.01*max((((2.191E4+(-2.115E9)*wrr))+(((-428.3)+4.045E7*wrr))*nfr)/nfr,1e-3)
+Rsub3_rf      =  Rsub2_rf
+Rdc_n33_rf    = max((86.7923*exp(-0.1713*wrr*1e6)),1e-3)
+Rsc_n33_rf    = max((86.7923*exp(-0.1713*wrr*1e6)),1e-3)
+Rds_rf	       = max(460.31*exp(-223066*wrr),1e-3)
+Djdb_AREA_rf  = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf    = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)                                                                                          
+Djsb_AREA_rf  = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf    = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)  
**********************************************
Lgate       ( 2 20) inductor  l=1p                        m=mrr
Rgate       (20 21) resistor  r=Rg_rf*(1+drg_n33_rf)      m=mrr
Cgd_ext     (21 11) capacitor c=Cgd_rf*(1+dcgdext_n33_rf) m=mrr
Cgs_ext     (21 31) capacitor c=Cgs_rf*(1+dcgsext_n33_rf) m=mrr
Cds_ext     (15 31) capacitor c=Cds_rf                    m=mrr
Rds         (11 15) resistor  r=Rds_rf                    m=mrr
Ldrain       (1 11) inductor  l=1p                        m=mrr
Lsource      (3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (12 11) ndio33_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (32 31) ndio33_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
djbdn  (4 5) diobpw_rf area=arpwr pj=pjpwr m=mrr
djpsub (6 5) dnwdio_rf area=ardnwr pj=pjdnwr m=mrr
**********************************************
Rsub1      (41  4)  resistor r=Rsub1_rf m=mrr
Rsub2      (41  12) resistor r=Rsub2_rf m=mrr
Rsub3      (41  32) resistor r=Rsub2_rf m=mrr
**********************************************
dnw33_6t_ckt_rf_r (11 21 31 41) n33_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model n33_ckt_r bsim4 type = n
**********************************************************************************************                                                                            
*                              3.3V CORE NMOS MODEL                               *                                                                            
**********************************************************************************************                                                                            
* GENERAL PARAMETERS                                                                                                                                           
*                                                                                                                                                              
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 0                 igbmod       = 0                 wpemod       = 0                 

***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 3.5e-007          lmax         = 0.0001            wmin         = 2.2e-007          
+wmax         = 0.0001            

***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               toxe         = 6.65e-009+dtoxe_n33_mismatch_rf         
+dtox         = 3.9e-010                                                          
+xj           = 1.6e-007          ndep         = 6.250661e+017     ngate        = 1.6e+020          
+rsh          = 12                

***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 1.02e-014         wln          = 1                 ww           = -2.677213e-015    
+wwn          = 1                 wwl          = -2.5e-021         ll           = -9.5e-015         
+lln          = 1                 lw           = 0                 lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 

***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-007         dwj          = 0                 
+xgw          = 0.31e-006                 xgl          = -1.38e-008                 
+xl           = -1.38e-008+dxl_n33_mismatch_rf                                                          
+xw           = 1.58e-008+dxw_n33_mismatch_rf                                                           

***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = 0.75619+dvth0_n33_mismatch_rf                                                           
+lvth0        = 2.0644e-009+dlvth0_n33_rf                                                      
+wvth0        = -1.6313e-008+dwvth0_n33_rf                                                     
+pvth0        = 2.393452e-015+dpvth0_n33_rf                                                    
+phin         = 0.15              k1           = 0.92              k2           = 0.0192267         
+lk2          = -1.7175e-008      wk2          = 1e-009            pk2          = 1.2125e-015       
+k3           = -1                lk3          = 3.247781e-006     wk3          = 1.174813e-006     
+pk3          = -2.895674e-013    k3b          = 2.7               lk3b         = -4.94e-006        
+wk3b         = 1.02e-006         pk3b         = 8.05e-013         w0           = 1.25e-006         
+lpe0         = 1.793508e-007     llpe0        = -3e-014           wlpe0        = -1.83375e-014     
+plpe0        = 2.8e-021          lpeb         = 0                 llpeb        = -1e-014           
+vbm          = -3                dvt0         = 1.977453          dvt1         = 0.81669           
+wdvt1        = 4.9e-009          dvt2         = -1.52658          dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            wint         = 3.409374e-008     lint         = 8.591858e-008     
+dwg          = -1e-009           wdwg         = 2.5e-016          dwb          = 0                 

***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.034389+du0_n33_mismatch_rf                                                            
+lu0          = -6.5037e-010+dlu0_n33_rf                                                       
+wu0          = 2.9719e-010+dwu0_n33_rf                                                        
+pu0          = 1.3e-016+dpu0_n33_rf                                                           
+ua           = -1.319673e-009    lua          = -3e-017           wua          = 4.255033e-017     
+pua          = -1.2e-023         ub           = 3.076021e-018     wub          = -1.578187e-025    
+pub          = 2e-033            uc           = 1.75496e-010      luc          = -6e-018           
+wuc          = -2e-017           puc          = -6e-025           ud           = 0                 
+eu           = 1.67              
+vsat         = 54975.69+dvsat_n33_mismatch_rf                                                          
+lvsat        = 0.0050622+dlvsat_n33_rf                                                        
+wvsat        = 0.001842913+dwvsat_n33_rf                                                      
+pvsat        = 1.370232e-010+dpvsat_n33_rf                                                    
+a0           = 1.446797          la0          = -3.3e-007         pa0          = 7e-014            
+ags          = 0.289501          lags         = 2.9e-007          wags         = -1.251297e-008    
+pags         = -1e-014           b0           = 8.604318e-008     lb0          = -6.913192e-014    
+wb0          = -4.812935e-014    pb0          = -1.044909e-020    b1           = 0                 
+lb1          = -1.606808e-014    wb1          = 1.713014e-013     pb1          = 8.347455e-021     
+keta         = -0.030075         lketa        = 1.391934e-009     pketa        = -7.784875e-015    
+a1           = 0                 a2           = 1                 

***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.147398+dvoff_n33_mismatch_rf         
+voffl        = -4.2e-009         minv         = -0.45             
+nfactor      = 1.066459          pnfactor     = -7e-015           eta0         = 0.08              
+etab         = -0.07             letab        = -1.7e-007         petab        = 2.5e-014          
+dsub         = 0.56              cit          = 4.634146e-005     cdsc         = 0.00024           
+cdscb        = 0                 cdscd        = 2e-005            

***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.26              pdiblc1      = 0.39              pdiblc2      = 0.000705          
+ppdiblc2     = -2.5e-017         pdiblcb      = 0                 drout        = 0.56              
+pscbe1       = 4.24e+008         pscbe2       = 1e-005            pvag         = 0                 
+delta        = 0                 ldelta       = 2e-009            fprout       = 0                 
+pdits        = 0                 pditsl       = 0                 pditsd       = 0                 

***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 549.89337         rdw          = 24                rdwmin       = 0                 
+rsw          = 24                rswmin       = 0                 prwg         = 0.108             
+prwb         = 0                 wr           = 1                 

***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 0                 alpha1       = 11.09775          lalpha1      = 2.123369e-005     
+beta0        = 25.056188         lbeta0       = 2e-006            

***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.002249          bigbacc      = 1.71e-007         cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0111            bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.00525           laigc        = -1.3e-010         waigc        = -1.2e-010         
+bigc         = 0.0003            cigc         = 0.075             dlcig        = 4e-009            
+aigsd        = 0.0045            waigsd       = -1e-010           bigsd        = 0.0001            
+cigsd        = 0.075             nigc         = 1                 poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 6.65e-009         

***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 0                 
+lagidl       = 0+dlagidl_n33_rf                                                               
+pagidl       = 0+dpagidl_n33_rf                                                               
+bgidl        = 2.3e+009          cgidl        = 0.5               egidl        = 0.8               

***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 6.25e+041         noib         = 5E+25        noic         = 8.75              
+em           = 4.1e+007          ef           = 1                 lintnoi      = 0                 
+ntnoi        = 1                 

***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_n33_rf)                     xrcrg1 = 10                       xrcrg2  = 8
+ngcon= 2
+rnoia = (max(0.01303+6.337*pwr(exp(10*(lrr*1e+6)),-0.8695)+0.56*pwr((wrr*1e+6),0.138),0.1))    tnoia = 0.1e+7    rnoib=0    tnoib=1.0e+7
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 1e-010+dcgdo_n33_rf                                                            
+cgso         = 1e-010+dcgso_n33_rf                                                            
+cgbo         = 0                 
+cgdl         = (2.6e-010+dcgdl_n33_rf)*0.8                                                          
+cgsl         = (2.6e-010+dcgsl_n33_rf)*0.8                                                          
+cf           = 7.55e-011+dcf_n33_rf
+clc          = 1e-007            cle          = 0.6               dlc          = 5.381e-008*(0.123*EXP(1404000*lr)+1)       
+dwc          = 0                 noff         = 2.2               lnoff        = 3.856e-007        
+voffcv       = -0.1184           lvoffcv      = -2.968e-008       acde         = 0.23814           
+moin         = 5.2               

***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.8              jss          = 4.1904e-007       jsws         = 3.9508e-013       
+jswgs        = 4.3285e-014       jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 
+jtsswgs      = 1.61e-009+djtsswgs_n33_rf                                                      
+jtsswgd      = 1.61e-009+djtsswgd_n33_rf                                                      
+njts         = 20                njtssw       = 20                njtsswg      = 20                
+xtss         = 0.02              xtsd         = 0.02              xtssws       = 0.02              
+xtsswd       = 0.02              xtsswgs      = 0.02              xtsswgd      = 0.02              
+vtss         = 10                vtsd         = 10                vtssws       = 10                
+vtsswd       = 10                vtsswgs      = 10                vtsswgd      = 10                
+tnjts        = 0               tnjtssw      = 0                 tnjtsswg     = 0                 
+cjs          = 0                                                        
+cjsws        = 0                                                      
+cjswgs       = 0                                                    
+mjs          = 0.32174           mjsws        = 0.0001727         mjswgs       = 0.36511           
+pbs          = 0.70384           pbsws        = 0.44462           pbswgs       = 0.59056           

***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.5              kt1          = -0.2565           
+lkt1         = 6e-009            pkt1         = 1.5e-015          kt2          = -0.0572           
+ua1          = 1e-009            ub1          = -1.29e-018        lub1         = -1e-025           
+wub1         = -1.17e-025        pub1         = 5e-032            uc1          = 5.6e-011          
+wuc1         = -1.68e-017        at           = 100000            lat          = -0.0157           
+pat          = 3e-010            njs          = 1.0296            xtis         = 3                 
+tpb          = 0.0016752         tpbsw        = 0.0009385         tpbswg       = 0.001502          
+tcj          = 0.00093975        tcjsw        = 0.00046393        tcjswg       = 0.0011153         
+tvoff        = 0.002             

***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 5.33e-006         sbref        = 5.33e-006         wlod         = 0                 
+ku0          = -2e-008           kvsat        = 1                 tku0         = 0                 
+lku0         = 5e-007            wku0         = 1e-006            pku0         = 0                 
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 6e-009            
+lkvth0       = 2e-007            wkvth0       = -5e-008           pkvth0       = 0                 
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                 

***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 1                 wec          = 1                 kvth0we      = 0            
+k2we         = 0                 ku0we        = 0           scref        = 1e-006            
*****************************************************************************************
* **
model ndio33_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
+dcap = 2 area = 4e-10 perim = 0.00008 tnom = 25 
+js = 4.1904e-007  isw = 3.9508e-013  expli = 1e+020 
+n = 1.0296  ns = 1.0296 rs = 2.8395e-010 jtun = 0 jtunsw = 0 
+ntun = 30 ibv = 2.50e+03 vb = 11.8 
+cj = 0.00086098+dcj_ndio33_rf cjsw = (9.677e-011+dcjsw_ndio33_rf)*0.5 vj = 0.70384 vjsw = 0.44462 
+fcs = 0 mj = 0.32174 mjsw = 0.16049 fc = 0 
+tt = 0 
+tlev = 1 tlevc = 1 tcv = 0 trs = 0.00065303 
+xti = 3 xtitun = 3 cta = 0.00093975 ctp = 0.00046393 
+pta = 0.0016752 ptp = 0.0009385 eg = 1.16 gap1 = 0.000702 
+gap2 = 1108 ttt1 = 0 ttt2 = 0 tm1 = 0 
+tm2 = 0 

model diobpw_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 1.0388e-006 isw = 1.4035e-013 vb = 15.5 ibv = 55.6 
+n = 1.1225 ns = 1.1225 rs = 1.8727e-010 
+cj = 0.00049858+dcj_diobpw_rf cjsw = 3.9867e-010+dcjsw_diobpw_rf vj = 0.67589 vjsw = 0.88873 
+fcs = 0 mj = 0.33041 mjsw = 0.444 fc = 0 
+tlev = 1 tlevc = 1 trs = 0.00035608 xti = 3 
+cta = 0.00090633 ctp = 0.00080455 pta = 0.001448 ptp = 0.0012196 
+eg = 1.16  tcv = -0.0005

model dnwdio_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-20
+area = 1.8e-008 perim = 0.00072 tnom = 25 
+js = 2.1632e-006 isw = 1.177e-012 vb = 16 ibv = 55.556 
+n = 1.0435 ns = 1.0435 rs = 1.3973e-007 
+cj = 0.00013824+dcj_dnwdio_rf cjsw = 4.1094e-010+dcjsw_dnwdio_rf vj = 0.52465 vjsw = 0.62598 
+fcs = 0 mj = 0.32294 mjsw = 0.35115 fc = 0 
+tlev = 1 tlevc = 1 trs = 1e-005 xti = 3 
+cta = 0.001326 ctp = 0.001221 pta = 0.0013127 ptp = 0.0015078 
+eg = 1.16 gap1 = 7.02e-04 tcv = -0.0006

ends dnw33_6t_ckt_rf_r


//* 3.3v pmos 
//* 1=drain,2=gate,3=source,4=bulk
inline subckt p33_ckt_rf_r (1 2 3 4)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.16u sbrr=1.16u sdrr=0.54u nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0 

**********************************************
+Cgd_rf = max(((0.9013*pwr(lrr*1e6,0.038)-0.8)*wrr*1e6+0.4911*pwr(lrr*1e6,0.1793))*nfr*1e-15,1e-18)
+Cgs_rf = max((0.4145*pwr(lrr*1e6,1.8456)+0.535)*nfr*(1.8232*pwr(nfr,-1.519)+0.987)*exp(wrr*1e6*(0.1426*pwr(nfr,-0.559)-0.01))*1e-15,1e-18)
+Cds_rf = max(1*((0.0306*pwr(lrr*1e6,-1.178)-0.03)*wrr*1e6-0.0143*lrr*1000000+0.0293)*nfr*1e-15,1e-18)
+Rg_rf  = max((195.55*pwr(nfr,-1.232)+4)*pwr(wrr*1000000,0.6293*pwr(nfr,-2.407)-0.306)*0.3205*pwr(lrr*1000000,-0.947),1e-3)
+Rsub1_rf = max(36.67*pwr(nfr,-0.252),1e-3)
+Rsub2_rf = max(94.041*exp(-0.036*nfr),1e-3)
+Djdb_AREA_rf = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf   = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)                                                                                          
+Djsb_AREA_rf = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf   = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)  
**********************************************
Lgate      (  2 20) inductor  l=1p                        m=mrr
Rgate      ( 20 21) resistor  r=Rg_rf*(1+drg_p33_rf)      m=mrr
Cgd_ext    ( 21 11) capacitor c=Cgd_rf*(1+dcgdext_p33_rf) m=mrr
Cgs_ext    ( 21 31) capacitor c=Cgs_rf*(1+dcgsext_p33_rf) m=mrr
Cds_ext    ( 15 31) capacitor c=Cds_rf                    m=mrr
Rds        ( 11 15) resistor  r=10                        m=mrr
Ldrain     (  1 11) inductor  l=1p                        m=mrr
Lsource    (  3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (11 12) pdio33_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (31 32) pdio33_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
**********************************************
Rsub1      (41  4 ) resistor  r= Rsub1_rf m=mrr
Rsub2      (41  12) resistor  r= Rsub2_rf m=mrr
Rsub3      (41  32) resistor  r= Rsub2_rf m=mrr
**********************************************
p33_ckt_rf_r (11 21 31 41) p33_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model p33_ckt_r bsim4 type = p

***********************************************************************************
*                             3.3V IO PMOS MODEL                                  *
***********************************************************************************
***********************************************************************************
*                             3.3V IO PMOS MODEL                                  *
***********************************************************************************
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 0                 igbmod       = 0                 wpemod       = 0                 
***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 3e-007            lmax         = 0.0001            wmin         = 2.2e-007          
+wmax         = 0.0001            
***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               toxe         = 6.64e-009+dtoxe_p33_rf_mismatch         
+dtox         = 1.7e-010                                                          
+xj           = 1.6e-007          ndep         = 1.6e+017          ngate        = 1e+020            
+rsh          = 12                
***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 0                 wln          = 1                 ww           = -1e-015           
+wwn          = 1                 wwl          = -1.61e-021        ll           = 1.258e-014        
+lln          = 1                 lw           = -4e-015           lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 
***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-7         dwj          = 0                 
+xgw          = 0.31e-6                 xgl          = -1.67e-008                 
+xl           = -1.67e-008+dxl_p33_rf_mismatch                                                          
+xw           = 1.58e-008+dxw_p33_rf_mismatch
+ngcon        = 2                                                          
***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = -0.69515+dvth0_p33_rf_mismatch                                                          
+lvth0        = 1.612e-007+dlvth0_p33_rf                                                       
+wvth0        = -3.1e-009+dwvth0_p33_rf                                                        
+pvth0        = 2.8e-015+dpvth0_p33_rf                                                         
+phin         = 0.11              k1           = 0.9               k2           = 0.042             
+lk2          = 4e-009            wk2          = -6e-009           k3           = 0.8               
+wk3          = 8.1e-007          pk3          = -9e-013           k3b          = 0.5               
+w0           = 2.839316e-006     lpe0         = 3.488847e-007     llpe0        = 7.382193e-015     
+plpe0        = 5.56e-022         lpeb         = -3e-008           llpeb        = -6e-015           
+plpeb        = 1e-022            vbm          = -3                dvt0         = 10                
+dvt1         = 0.5               dvt2         = -0.002            dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            wint         = 2e-008            lint         = -4.35e-008        
+dwg          = 0                 wdwg         = 1e-016            pdwg         = 1.4e-022          
+dwb          = 0                 
***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.011408+du0_p33_rf_mismatch                                                            
+lu0          = -1.3e-010+dlu0_p33_rf                                                          
+wu0          = 4.6465e-010+dwu0_p33_rf                                                        
+pu0          = -2.44e-016+dpu0_p33_rf                                                         
+ua           = 9.421845e-010     lua          = -2.346753e-016    wua          = -6e-017           
+pua          = -4.25e-023        ub           = 8.107345e-019     lub          = 4.237495e-025     
+wub          = -1.53e-025        pub          = -5e-033           uc           = -3.125e-011       
+luc          = 5.845e-017        wuc          = -2.0625e-017      puc          = -1.68e-024        
+ud           = 0                 eu           = 1                 
+vsat         = 71203.72+dvsat_p33_rf_mismatch                                                          
+lvsat        = 0.0131721+dlvsat_p33_rf                                                        
+wvsat        = -0.001+dwvsat_p33_rf                                                           
+pvsat        = -1.17e-009+dpvsat_p33_rf                                                       
+a0           = 1.1               la0          = 5e-008            ags          = 0.14              
+lags         = 2e-007            wags         = -1.3e-008         b0           = -1e-008           
+wb0          = 1e-015            b1           = 0                 keta         = -0.004635593      
+lketa        = -1.5e-008         wketa        = 3.194915e-009     pketa        = 4.1e-016          
+a1           = 0.05              la1          = -2.5e-008         pa1          = -3e-015           
+a2           = 1                 
***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.153+dvoff_p33_rf_mismatch            pvoff        = 1e-015            voffl        = 2.411908e-008     
+minv         = -0.0971895        lminv        = 2e-007            wminv        = -1e-007           
+pminv        = 2.915685e-014     nfactor      = 0.357             lnfactor     = -4.256665e-008    
+wnfactor     = 2.1e-007          pnfactor     = -5.6e-014         eta0         = 0.0001+deta0_p33_rf_mismatch            
+leta0        = 3.1e-008          peta0        = 2e-015            etab         = -0.113            
+petab        = -1.2e-014         dsub         = 0.56              cit          = 0.00155           
+lcit         = 2e-010            cdsc         = 0.00024           cdscb        = 0                 
+cdscd        = 2e-005            
***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.65              lpclm        = -5.75e-008        ppclm        = 4.8e-015          
+pdiblc1      = 0.07              pdiblc2      = 0.0001            lpdiblc2     = -2e-011           
+wpdiblc2     = 5e-011            ppdiblc2     = 1.2e-016          pdiblcb      = 0                 
+drout        = 0.56              pscbe1       = 4.24e+008         pscbe2       = 1e-010            
+pvag         = 0                 delta        = 0.01              ldelta       = 3e-009            
+fprout       = 0                 pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 
***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 1300              prdsw        = -5e-011           rdw          = 24                
+rdwmin       = 0                 rsw          = 24                rswmin       = 0                 
+prwg         = 1                 prwb         = 0                 wr           = 1                 
***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 0.0044            alpha1       = 156.4             lalpha1      = -0.0044394        
+walpha1      = 0.000117          palpha1      = -3.37e-011        beta0        = 40.085            
+lbeta0       = -3.2e-006         wbeta0       = 1.4e-006          
***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.003             bigbacc      = 1.71e-007         cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0111            bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.0034            laigc        = -1e-010           waigc        = -8e-011           
+paigc        = -3e-018           bigc         = 0.00011           lbigc        = -3e-012           
+cigc         = 0.048             lcigc        = -1e-009           dlcig        = 4e-009            
+aigsd        = 0.0032            laigsd       = -1.38e-010        waigsd       = -9e-011           
+paigsd       = 1.3e-017          bigsd        = 0.0001            lbigsd       = 5e-011            
+wbigsd       = 2e-011            pbigsd       = -2e-018           cigsd        = 0.03              
+lcigsd       = 4.3e-008          nigc         = 2                 poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 6.64e-009         
***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 7.5828e-013+dagidl_p33_rf                                                      
+lagidl       = 3e-019+dlagidl_p33_rf                                                          
+wagidl       = 9e-019+dwagidl_p33_rf                                                          
+pagidl       = -2e-025+dpagidl_p33_rf                                                         
+bgidl        = 8.8e+008          cgidl        = 2                 egidl        = 0.63              
***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 3.156e+041        noib         = 3.1875e+024       noic         = 8e+009            
+em           = 3.075e+007        ef           = 1.1               lintnoi      = 0                 
+ntnoi        = 1                 
***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_p33_rf)                     xrcrg1 =8             xrcrg2  = 9
+rnoia = (max(0.224+7.855*pwr(exp(10*(lrr*1e+6)),-1.445)+0.309*pwr((wrr*1e+6),0.041),0.1))    tnoia = 1.3e+7    rnoib=0    tnoib=1.0e+7      
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 1e-010+dcgdo_p33_rf                                                            
+cgso         = 1e-010+dcgso_p33_rf                                                            
+cgbo         = 0                 
+cgdl         = 2.52e-010*0.8+dcgdl_p33_rf                                                         
+cgsl         = 2.52e-010*0.8+dcgsl_p33_rf                                                         
+cf           = 3.05e-011+dcf_p33_rf                                                           
+clc          = 0           cle          = 0.6               dlc          = 5.2375e-008*1       
+dwc          = 0                 noff         = 2             lnoff        = 2.31e-007
+voffcv       = -0.01             lvoffcv      = -1.575e-008       acde         = 0.37             
+moin         = 5.2  
*
***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.3              jss          = 1.06e-007         jsws         = 4.97e-014         
+jswgs        = 1.08e-014         jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 7e-011            
+jtsswgd      = 7e-011            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              vtss         = 10                vtsd         = 10                
+vtssws       = 10                vtsswd       = 10                vtsswgs      = 10                
+vtsswgd      = 10                tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                 
+cjs          = 0                                                           
+cjsws        = 0                                                        
+cjswgs       = 0                                                     
+mjs          = 0.398             mjsws        = 0.30364           mjswgs       = 0.32993           
+pbs          = 0.82134           pbsws        = 0.63646           pbswgs       = 0.56135           
***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.3              kt1          = -0.33  
+wkt1         = -6E-9                        
+lkt1         = -1e-008           kt2          = -0.046            lkt2         = 5e-009            
+ua1          = -1e-025           ub1          = -1.8e-018         lub1         = -6e-026           
+wub1         = 2e-025            pub1         = 1.2e-032          uc1          = -5.04e-011        
+luc1         = -4.1e-017         wuc1         = 2.6e-017          puc1         = -2e-024           
+at           = 100000            lat          = -0.028            wat          = 0.0098            
+pat          = -8e-009           njs          = 0.99891           xtis         = 3                 
+tpb          = 0.0015412         tpbsw        = 0.0022178         tpbswg       = 0.0013894         
+tcj          = 0.00092673        tcjsw        = 0.0012244         tcjswg       = 0.00084165        
***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 5.33e-006         sbref        = 5.33e-006         wlod         = 0                 
+ku0          = 8.1e-008          kvsat        = 1                 tku0         = 0                 
+lku0         = 2.8e-007          wku0         = -7e-008           pku0         = -1.2e-014         
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 1e-009            
+lkvth0       = 2.9e-007          wkvth0       = 5e-006            pkvth0       = 0                 
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                 
***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 1                 wec          = 1                 kvth0we      = 0            
+k2we         = 0                 ku0we        = 0           scref        = 1e-006 

***********************  

model pdio33_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 4e-010 perim = 8e-005 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 1.0586e-007 isw = 4.9737e-014 vb = 11.0 ibv = 2500 
+n = 0.99891 ns = 0.99891 rs = 5.87e-010 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = 0.001044+dcjs_p33_rf cjp = 8.5736e-011+dcjsws_p33_rf vj = 0.82134 vjsw = 0.63646 
+fcs = 0 mj = 0.398 mjsw = 0.30364 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 tcv = 0 trs = 0.002833 
+xti = 3 cta = 0.00092673 ctp = 0.0012244 pta = 0.0015412 
+ptp = 0.0022178 eg = 1.16 

ends p33_ckt_rf_r

//* 3.3v pmos 
//* 1=drain,2=gate,3=source,4=bulk,5=psub
inline subckt p33_5t_ckt_rf_r (1 2 3 4 5)
parameters wrr=1e-6 lrr=1e-6 nfr=1 sarr=1.16u sbrr=1.16u sdrr=0.54u nrdrr=0.001 nrsrr=0.001 mrr=1 scarr=0 scbrr=0 sccrr=0  arnwr=1e-12 pjnwr=4e-6

**********************************************
+Cgd_rf = max(((0.9013*pwr(lrr*1e6,0.038)-0.8)*wrr*1e6+0.4911*pwr(lrr*1e6,0.1793))*nfr*1e-15,1e-18)
+Cgs_rf = max((0.4145*pwr(lrr*1e6,1.8456)+0.535)*nfr*(1.8232*pwr(nfr,-1.519)+0.987)*exp(wrr*1e6*(0.1426*pwr(nfr,-0.559)-0.01))*1e-15,1e-18)
+Cds_rf = max(1*((0.0306*pwr(lrr*1e6,-1.178)-0.03)*wrr*1e6-0.0143*lrr*1000000+0.0293)*nfr*1e-15,1e-18)
+Rg_rf  = max((195.55*pwr(nfr,-1.232)+4)*pwr(wrr*1000000,0.6293*pwr(nfr,-2.407)-0.306)*0.3205*pwr(lrr*1000000,-0.947),1e-3)
+Rsub1_rf = max(36.67*pwr(nfr,-0.252),1e-3)
+Rsub2_rf = max(94.041*exp(-0.036*nfr),1e-3)
+Djdb_AREA_rf = int(0.5*(nfr+1))*(wrr*(0.54-2*0.07)*1e-6)                                                                                                      
+Djdb_PJ_rf   = int(0.5*(nfr+1))*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)                                                                                          
+Djsb_AREA_rf = int(0.5*nfr+1)*wrr*(0.54-2*0.07)*1e-6                                                                                                          
+Djsb_PJ_rf   = int(0.5*nfr+1)*(2*(0.54-2*0.07)*1e-6+2*wrr*4.71)  
**********************************************
Lgate      (  2 20) inductor  l=1p                        m=mrr
Rgate      ( 20 21) resistor  r=Rg_rf*(1+drg_p33_rf)      m=mrr
Cgd_ext    ( 21 11) capacitor c=Cgd_rf*(1+dcgdext_p33_rf) m=mrr
Cgs_ext    ( 21 31) capacitor c=Cgs_rf*(1+dcgsext_p33_rf) m=mrr
Cds_ext    ( 15 31) capacitor c=Cds_rf                    m=mrr
Rds        ( 11 15) resistor  r=10                        m=mrr
Ldrain     (  1 11) inductor  l=1p                        m=mrr
Lsource    (  3 31) inductor  l=1p                        m=mrr
**********************************************
Djdb  (11 12) pdio33_rf AREA=Djdb_AREA_rf PJ=Djdb_PJ_rf m=mrr
Djsb  (31 32) pdio33_rf AREA=Djsb_AREA_rf PJ=Djsb_PJ_rf m=mrr
Djnw  (5 4  ) nwdio_rf  AREA=arnwr PJ=pjnwr               m=mrr 
**********************************************
Rsub1      (41  4 ) resistor  r= Rsub1_rf m=mrr
Rsub2      (41  12) resistor  r= Rsub2_rf m=mrr
Rsub3      (41  32) resistor  r= Rsub2_rf m=mrr
**********************************************
p33_5t_ckt_rf_r (11 21 31 41) p33_ckt_r w=(wrr*nfr) l=lrr sa=sarr sb=sbrr sd=sdrr as=0 ad=0 ps=0 pd=0 nrd=nrdrr nrs=nrsrr sca=scarr scb=scbrr scc=sccrr nf=nfr m=mrr
model p33_ckt_r bsim4 type = p

***********************************************************************************
*                             3.3V IO PMOS MODEL                                  *
***********************************************************************************
***************************************************************************
*             Model Selector Parameter
***************************************************************************
+level        = 54                version      = 4.5               binunit      = 2                 
+paramchk     = 1                 mobmod       = 0                 capmod       = 2                 
+rgatemod     = 3                 geomod       = 0                 rgeomod      = 1                 
+diomod       = 2                 rdsmod       = 0                 rbodymod     = 0                 
+fnoimod      = 1                 tnoimod      = 1                 tempmod      = 0                 
+permod       = 1                 acnqsmod     = 0                 trnqsmod     = 0                 
+igcmod       = 0                 igbmod       = 0                 wpemod       = 0                 
***************************************************************************
*             Geometry Range Parameter
***************************************************************************
+lmin         = 3e-007            lmax         = 0.0001            wmin         = 2.2e-007          
+wmax         = 0.0001            
***************************************************************************
*             Process Parameter
***************************************************************************
+epsrox       = 3.9               toxe         = 6.64e-009+dtoxe_p33_rf_mismatch         
+dtox         = 1.7e-010                                                          
+xj           = 1.6e-007          ndep         = 1.6e+017          ngate        = 1e+020            
+rsh          = 12                
***************************************************************************
*             dW and dL Parameter
***************************************************************************
+wl           = 0                 wln          = 1                 ww           = -1e-015           
+wwn          = 1                 wwl          = -1.61e-021        ll           = 1.258e-014        
+lln          = 1                 lw           = -4e-015           lwn          = 1                 
+lwl          = 0                 llc          = 0                 lwc          = 0                 
+lwlc         = 0                 wlc          = 0                 wwc          = 0                 
+wwlc         = 0                 
***************************************************************************
*             Layout-Dependent Parasitics Model Parameter
***************************************************************************
+dmcg         = 2.7e-007          dmci         = 2.7e-7         dwj          = 0                 
+xgw          = 0.31e-6                 xgl          = -1.67e-008                 
+xl           = -1.67e-008+dxl_p33_rf_mismatch                                                          
+xw           = 1.58e-008+dxw_p33_rf_mismatch
+ngcon        = 2                                                          
***************************************************************************
*             BASIC: Vth Related  Parameter
***************************************************************************
+vth0         = -0.69515+dvth0_p33_rf_mismatch                                                          
+lvth0        = 1.612e-007+dlvth0_p33_rf                                                       
+wvth0        = -3.1e-009+dwvth0_p33_rf                                                        
+pvth0        = 2.8e-015+dpvth0_p33_rf                                                         
+phin         = 0.11              k1           = 0.9               k2           = 0.042             
+lk2          = 4e-009            wk2          = -6e-009           k3           = 0.8               
+wk3          = 8.1e-007          pk3          = -9e-013           k3b          = 0.5               
+w0           = 2.839316e-006     lpe0         = 3.488847e-007     llpe0        = 7.382193e-015     
+plpe0        = 5.56e-022         lpeb         = -3e-008           llpeb        = -6e-015           
+plpeb        = 1e-022            vbm          = -3                dvt0         = 10                
+dvt1         = 0.5               dvt2         = -0.002            dvtp0        = 0                 
+dvtp1        = 0                 dvt0w        = 0                 dvt1w        = 5300000           
+dvt2w        = -0.032            wint         = 2e-008            lint         = -4.35e-008        
+dwg          = 0                 wdwg         = 1e-016            pdwg         = 1.4e-022          
+dwb          = 0                 
***************************************************************************
*             BASIC: Mobility Related Parameter
***************************************************************************
+u0           = 0.011408+du0_p33_rf_mismatch                                                            
+lu0          = -1.3e-010+dlu0_p33_rf                                                          
+wu0          = 4.6465e-010+dwu0_p33_rf                                                        
+pu0          = -2.44e-016+dpu0_p33_rf                                                         
+ua           = 9.421845e-010     lua          = -2.346753e-016    wua          = -6e-017           
+pua          = -4.25e-023        ub           = 8.107345e-019     lub          = 4.237495e-025     
+wub          = -1.53e-025        pub          = -5e-033           uc           = -3.125e-011       
+luc          = 5.845e-017        wuc          = -2.0625e-017      puc          = -1.68e-024        
+ud           = 0                 eu           = 1                 
+vsat         = 71203.72+dvsat_p33_rf_mismatch                                                          
+lvsat        = 0.0131721+dlvsat_p33_rf                                                        
+wvsat        = -0.001+dwvsat_p33_rf                                                           
+pvsat        = -1.17e-009+dpvsat_p33_rf                                                       
+a0           = 1.1               la0          = 5e-008            ags          = 0.14              
+lags         = 2e-007            wags         = -1.3e-008         b0           = -1e-008           
+wb0          = 1e-015            b1           = 0                 keta         = -0.004635593      
+lketa        = -1.5e-008         wketa        = 3.194915e-009     pketa        = 4.1e-016          
+a1           = 0.05              la1          = -2.5e-008         pa1          = -3e-015           
+a2           = 1                 
***************************************************************************
*             BASIC: Subthreshold Related Parameter
***************************************************************************
+voff         = -0.153+dvoff_p33_rf_mismatch            pvoff        = 1e-015            voffl        = 2.411908e-008     
+minv         = -0.0971895        lminv        = 2e-007            wminv        = -1e-007           
+pminv        = 2.915685e-014     nfactor      = 0.357             lnfactor     = -4.256665e-008    
+wnfactor     = 2.1e-007          pnfactor     = -5.6e-014         eta0         = 0.0001+deta0_p33_rf_mismatch            
+leta0        = 3.1e-008          peta0        = 2e-015            etab         = -0.113            
+petab        = -1.2e-014         dsub         = 0.56              cit          = 0.00155           
+lcit         = 2e-010            cdsc         = 0.00024           cdscb        = 0                 
+cdscd        = 2e-005            
***************************************************************************
*             BASIC: Output Resistance Related Parameter
***************************************************************************
+pclm         = 0.65              lpclm        = -5.75e-008        ppclm        = 4.8e-015          
+pdiblc1      = 0.07              pdiblc2      = 0.0001            lpdiblc2     = -2e-011           
+wpdiblc2     = 5e-011            ppdiblc2     = 1.2e-016          pdiblcb      = 0                 
+drout        = 0.56              pscbe1       = 4.24e+008         pscbe2       = 1e-010            
+pvag         = 0                 delta        = 0.01              ldelta       = 3e-009            
+fprout       = 0                 pdits        = 0                 pditsl       = 0                 
+pditsd       = 0                 
***************************************************************************
*             Asymmetric and Bias-Dependent
***************************************************************************
+rdsw         = 1300              prdsw        = -5e-011           rdw          = 24                
+rdwmin       = 0                 rsw          = 24                rswmin       = 0                 
+prwg         = 1                 prwb         = 0                 wr           = 1                 
***************************************************************************
*             Impact Ionization Current Model Parameters
***************************************************************************
+alpha0       = 0.0044            alpha1       = 156.4             lalpha1      = -0.0044394        
+walpha1      = 0.000117          palpha1      = -3.37e-011        beta0        = 40.085            
+lbeta0       = -3.2e-006         wbeta0       = 1.4e-006          
***************************************************************************
*             Gate Dielectric Tunneling Current
***************************************************************************
+aigbacc      = 0.003             bigbacc      = 1.71e-007         cigbacc      = 0.075             
+nigbacc      = 1                 aigbinv      = 0.0111            bigbinv      = 0.000949          
+cigbinv      = 0.006             eigbinv      = 1.1               nigbinv      = 3                 
+aigc         = 0.0034            laigc        = -1e-010           waigc        = -8e-011           
+paigc        = -3e-018           bigc         = 0.00011           lbigc        = -3e-012           
+cigc         = 0.048             lcigc        = -1e-009           dlcig        = 4e-009            
+aigsd        = 0.0032            laigsd       = -1.38e-010        waigsd       = -9e-011           
+paigsd       = 1.3e-017          bigsd        = 0.0001            lbigsd       = 5e-011            
+wbigsd       = 2e-011            pbigsd       = -2e-018           cigsd        = 0.03              
+lcigsd       = 4.3e-008          nigc         = 2                 poxedge      = 1                 
+pigcd        = 1                 ntox         = 1                 toxref       = 6.64e-009         
***************************************************************************
*             GIDL Effect Parameters
***************************************************************************
+agidl        = 7.5828e-013+dagidl_p33_rf                                                      
+lagidl       = 3e-019+dlagidl_p33_rf                                                          
+wagidl       = 9e-019+dwagidl_p33_rf                                                          
+pagidl       = -2e-025+dpagidl_p33_rf                                                         
+bgidl        = 8.8e+008          cgidl        = 2                 egidl        = 0.63              
***************************************************************************
*             Flicker Noise Model Parameter
***************************************************************************
+noia         = 3.156e+041        noib         = 3.1875e+024       noic         = 8e+009            
+em           = 3.075e+007        ef           = 1.1               lintnoi      = 0                 
+ntnoi        = 1                 
***************************************************************************
*             High-Speed RF Model Parameters
***************************************************************************
+rshg = (rshg_p33_rf)                     xrcrg1 =8             xrcrg2  = 9
+rnoia = (max(0.224+7.855*pwr(exp(10*(lrr*1e+6)),-1.445)+0.309*pwr((wrr*1e+6),0.041),0.1))    tnoia = 1.3e+7    rnoib=0    tnoib=1.0e+7      
***************************************************************************
*             Capacitance Parameter
***************************************************************************
+xpart        = 0                 
+cgdo         = 1e-010+dcgdo_p33_rf                                                            
+cgso         = 1e-010+dcgso_p33_rf                                                            
+cgbo         = 0                 
+cgdl         = 2.52e-010*0.8+dcgdl_p33_rf                                                         
+cgsl         = 2.52e-010*0.8+dcgsl_p33_rf                                                         
+cf           = 3.05e-011+dcf_p33_rf                                                           
+clc          = 0           cle          = 0.6               dlc          = 5.2375e-008*1       
+dwc          = 0                 noff         = 2             lnoff        = 2.31e-007
+voffcv       = -0.01             lvoffcv      = -1.575e-008       acde         = 0.37             
+moin         = 5.2  
*
***************************************************************************
*             Souce|Drain Junction Diode Model Parameter
***************************************************************************
+ijthsrev     = 0.1               ijthsfwd     = 0.1               xjbvs        = 1                 
+bvs          = 11.3              jss          = 1.06e-007         jsws         = 4.97e-014         
+jswgs        = 1.08e-014         jtss         = 0                 jtsd         = 0                 
+jtssws       = 0                 jtsswd       = 0                 jtsswgs      = 7e-011            
+jtsswgd      = 7e-011            njts         = 20                njtssw       = 20                
+njtsswg      = 20                xtss         = 0.02              xtsd         = 0.02              
+xtssws       = 0.02              xtsswd       = 0.02              xtsswgs      = 0.02              
+xtsswgd      = 0.02              vtss         = 10                vtsd         = 10                
+vtssws       = 10                vtsswd       = 10                vtsswgs      = 10                
+vtsswgd      = 10                tnjts        = 0                 tnjtssw      = 0                 
+tnjtsswg     = 0                 
+cjs          = 0                                                           
+cjsws        = 0                                                        
+cjswgs       = 0                                                     
+mjs          = 0.398             mjsws        = 0.30364           mjswgs       = 0.32993           
+pbs          = 0.82134           pbsws        = 0.63646           pbswgs       = 0.56135           
***************************************************************************
*             Temperature coefficient
***************************************************************************
+tnom         = 25                ute          = -1.3              kt1          = -0.33  
+wkt1         = -6E-9                        
+lkt1         = -1e-008           kt2          = -0.046            lkt2         = 5e-009            
+ua1          = -1e-025           ub1          = -1.8e-018         lub1         = -6e-026           
+wub1         = 2e-025            pub1         = 1.2e-032          uc1          = -5.04e-011        
+luc1         = -4.1e-017         wuc1         = 2.6e-017          puc1         = -2e-024           
+at           = 100000            lat          = -0.028            wat          = 0.0098            
+pat          = -8e-009           njs          = 0.99891           xtis         = 3                 
+tpb          = 0.0015412         tpbsw        = 0.0022178         tpbswg       = 0.0013894         
+tcj          = 0.00092673        tcjsw        = 0.0012244         tcjswg       = 0.00084165        
***************************************************************************
*             Stress Effect Related Parameter
***************************************************************************
+saref        = 5.33e-006         sbref        = 5.33e-006         wlod         = 0                 
+ku0          = 8.1e-008          kvsat        = 1                 tku0         = 0                 
+lku0         = 2.8e-007          wku0         = -7e-008           pku0         = -1.2e-014         
+llodku0      = 1                 wlodku0      = 1                 kvth0        = 1e-009            
+lkvth0       = 2.9e-007          wkvth0       = 5e-006            pkvth0       = 0                 
+llodvth      = 1                 wlodvth      = 1                 stk2         = 0                 
+lodk2        = 1                 steta0       = 0                 lodeta0      = 1                 
***************************************************************************
*             Well Proximity Effect Model Parameters
***************************************************************************
+web          = 1                 wec          = 1                 kvth0we      = 0            
+k2we         = 0                 ku0we        = 0           scref        = 1e-006 

***********************  

model pdio33_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 4e-010 perim = 8e-005 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 1.0586e-007 isw = 4.9737e-014 vb = 11.0 ibv = 2500 
+n = 0.99891 ns = 0.99891 rs = 5.87e-010 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = 0.001044+dcjs_p33_rf cjp = 8.5736e-011+dcjsws_p33_rf vj = 0.82134 vjsw = 0.63646 
+fcs = 0 mj = 0.398 mjsw = 0.30364 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 tcv = 0 trs = 0.002833 
+xti = 3 cta = 0.00092673 ctp = 0.0012244 pta = 0.0015412 
+ptp = 0.0022178 eg = 1.16 

// **  
model nwdio_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 9.6e-009 perim = 4e-004 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 2.3733e-006 isw = 2.9142e-014 vb = 15 ibv = 104 
+n = 1.085 ns = 1.085 rs = 8.4602e-009 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = 0.000131+dcj_nwdio_rf cjp = 5.0047e-010+dcjp_nwdio_rf vj = 0.41624 vjsw = 0.81575 
+fcs = 0 mj = 0.26295 mjsw = 0.377 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 trs = 0.0004 xti = 3 
+cta = 0.0017608 ctp = 0.0012659 pta = 0.00155 ptp = 0.0022128 
+eg = 1.16 
// *
//
ends p33_5t_ckt_rf_r

