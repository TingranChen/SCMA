//* 
//* No part of this file can be released without the consent of SMIC.                                                                                                                                                                                            
//*                                                                                                                                                                                                                                                              
//************************************************************************************************************                                                                                                                                                   
//* smic 0.18um mixed signal 1p6m 1.8v/3.3v spice model(for SPECTRE only) //*                                                                                                                                                     
//************************************************************************************************************                                                                                                                                                   
//*                                                                                                                                                                                                                                                              
//* Release version    : 1.11                                                                                                                                                                                                                                     
//*                                                                                                                                                                                                                                                              
//* Release date       : 17/03/2015                                                                                                                                                                                                                              
//*                                                                                                                                                                                                                                                              
//* Simulation tool    : Cadence spectre V6.1.1.399                                                                                                                                                                                                 
//*                                                                                                                                                                                                                                                              
//*  Inductor   :                                                                                                                                                                                                                                                
//* *  *------------------------*---------------------------------------------------------*
//*    |  Turn, Radius & Width  |  T=2~7.5 step 0.5,W=3~15um,R=1.7071*W+11.878~90um       |
//* *  *------------------------*---------------------------------------------------------*
//*    |        Model Name      |           ind_rf_psub                                  |            
//* *  *------------------------*---------------------------------------------------------*
simulator lang=spectre  insensitive=yes
subckt ind_rf_psub (PLUS MINUS PSUB)
parameters R=6e-05 radius_=0.0111111*(R/1e-06-0) w=8e-06 w_=0.0666667*(w/1e-06-0) n=3  \
T0=(n==2.5) \
T1=(radius_>=0.444722) \
T2=(w_+6.944444e-01*radius_>=0.909235) \
T3=(w_>=0.6004) \
T4=(radius_>=0.444167) \
T5=(radius_>=0.7225) \
T6=(w_+6.944444e-01*radius_>=0.908049) \
T7=(w_>=0.5996) \
T8=(radius_>=0.721944) \
T9=(n==2) \
T10=(n==3.5) \
T11=(n==3) \
T12=(n==4.5) \
T13=(n==4) \
T14=(n==5.5) \
T15=(n==5) \
T16=(n==6.5) \
T17=(n==6) \
T18=(n==7.5) \
T19=(n==7) \
S0=T0*(1-T1)*(1-T2) \
noS0=(1-S0) \
S1=T0*(1-T3)*T4*(1-T5)*noS0 \
noS1=(1-S1)*noS0 \
S2=T0*T6*T7*(1-T5)*noS1 \
noS2=(1-S2)*noS1 \
S3=T0*(1-T3)*T8*noS2 \
noS3=(1-S3)*noS2 \
S4=T0*T8*T7*noS3 \
noS4=(1-S4)*noS3 \
S5=T9*(1-T1)*(1-T2)*noS4 \
noS5=(1-S5)*noS4 \
S6=T9*(1-T3)*T4*(1-T5)*noS5 \
noS6=(1-S6)*noS5 \
S7=T9*T6*T7*(1-T5)*noS6 \
noS7=(1-S7)*noS6 \
S8=T9*(1-T3)*T8*noS7 \
noS8=(1-S8)*noS7 \
S9=T9*T8*T7*noS8 \
noS9=(1-S9)*noS8 \
S10=T10*(1-T1)*noS9 \
noS10=(1-S10)*noS9 \
S11=T10*T4*(1-T5)*noS10 \
noS11=(1-S11)*noS10 \
S12=T10*T8*noS11 \
noS12=(1-S12)*noS11 \
S13=T11*(1-T1)*(1-T2)*noS12 \
noS13=(1-S13)*noS12 \
S14=T11*(1-T3)*T4*(1-T5)*noS13 \
noS14=(1-S14)*noS13 \
S15=T11*T6*T7*(1-T5)*noS14 \
noS15=(1-S15)*noS14 \
S16=T11*(1-T3)*T8*noS15 \
noS16=(1-S16)*noS15 \
S17=T11*T8*T7*noS16 \
noS17=(1-S17)*noS16 \
S18=T12*(1-T1)*noS17 \
noS18=(1-S18)*noS17 \
S19=T12*T4*(1-T5)*noS18 \
noS19=(1-S19)*noS18 \
S20=T12*T8*noS19 \
noS20=(1-S20)*noS19 \
S21=T13*(1-T1)*noS20 \
noS21=(1-S21)*noS20 \
S22=T13*T4*(1-T5)*noS21 \
noS22=(1-S22)*noS21 \
S23=T13*T8*noS22 \
noS23=(1-S23)*noS22 \
S24=T14*(1-T1)*noS23 \
noS24=(1-S24)*noS23 \
S25=T14*T4*(1-T5)*noS24 \
noS25=(1-S25)*noS24 \
S26=T14*T8*noS25 \
noS26=(1-S26)*noS25 \
S27=T15*(1-T1)*noS26 \
noS27=(1-S27)*noS26 \
S28=T15*T4*(1-T5)*noS27 \
noS28=(1-S28)*noS27 \
S29=T15*T8*noS28 \
noS29=(1-S29)*noS28 \
S30=T16*(1-T1)*noS29 \
noS30=(1-S30)*noS29 \
S31=T16*T4*(1-T5)*noS30 \
noS31=(1-S31)*noS30 \
S32=T16*T8*noS31 \
noS32=(1-S32)*noS31 \
S33=T17*(1-T1)*noS32 \
noS33=(1-S33)*noS32 \
S34=T17*T4*(1-T5)*noS33 \
noS34=(1-S34)*noS33 \
S35=T17*T8*noS34 \
noS35=(1-S35)*noS34 \
S36=T18*(1-T1)*noS35 \
noS36=(1-S36)*noS35 \
S37=T18*T4*(1-T5)*noS36 \
noS37=(1-S37)*noS36 \
S38=T18*T8*noS37 \
noS38=(1-S38)*noS37 \
S39=T19*(1-T1)*noS38 \
noS39=(1-S39)*noS38 \
S40=T19*T4*(1-T5)*noS39 \
noS40=(1-S40)*noS39 \
S41=T19*T8*noS40 \
noS41=(1-S41)*noS40 \
V0_part1=3.985390e-01*S0+(-2.288517e+00)*S1+5.634825e-01*S2+(-1.958793e+00)*S3+(-5.865080e+00)*S4+3.437324e+00*S5+(-1.574767e-01)*S6+1.802128e+00*S7+(-5.730958e-01)*S8+(-7.648988e+00)*S9 \
V0_part2=V0_part1+1.617362e+00*S10+0.000000e+00*S11+(-3.488074e+00)*S12+(-3.088809e-01)*S13+2.983931e+00*S14+(-9.590618e-01)*S15+0.000000e+00*S16+(-3.676782e+00)*S17+0.000000e+00*S18+0.000000e+00*S19 \
V0_part3=V0_part2+(-2.627158e+00)*S20+0.000000e+00*S21+(-2.150748e+00)*S22+0.000000e+00*S23+(-9.755381e-01)*S24+(-3.022077e+00)*S25+0.000000e+00*S26+0.000000e+00*S27+(-1.582405e-01)*S28+4.029592e-02*S29 \
V0_part4=V0_part3+(-1.436199e+00)*S30+(-1.148209e-01)*S31+0.000000e+00*S32+(-7.222603e-02)*S33+1.430872e-02*S34+(-1.801973e-01)*S35+0.000000e+00*S36+0.000000e+00*S37+(-3.739412e+00)*S38+1.262085e+00*S39 \
V0=V0_part4+0.000000e+00*S40+(-1.076697e+01)*S41 \
V1_part1=7.658523e+00*S0+1.964781e+01*S1+5.573710e+00*S2+6.015491e+00*S3+2.101111e+01*S4+3.010454e+00*S5+1.771942e+01*S6+3.395943e+00*S7+1.758692e+01*S8+2.201347e+01*S9 \
V1_part2=V1_part1+1.094204e+00*S10+0.000000e+00*S11+1.826252e+01*S12+5.215191e+00*S13+2.247533e-03*S14+1.591490e+01*S15+0.000000e+00*S16+2.091132e+01*S17+0.000000e+00*S18+0.000000e+00*S19 \
V1_part3=V1_part2+1.218216e+01*S20+0.000000e+00*S21+1.648662e+01*S22+0.000000e+00*S23+2.020181e+01*S24+1.912790e+01*S25+0.000000e+00*S26+0.000000e+00*S27+1.050529e+01*S28+4.731693e+00*S29 \
V1_part4=V1_part3+1.656252e+01*S30+7.519784e-02*S31+0.000000e+00*S32+1.520140e+01*S33+1.527080e+01*S34+1.444997e+01*S35+0.000000e+00*S36+0.000000e+00*S37+1.588514e+01*S38+1.366808e+01*S39 \
V1=V1_part4+0.000000e+00*S40+1.513587e+01*S41 \
V2_part1=3.162898e-01*S0+4.493995e+00*S1+2.816422e+00*S2+4.989757e+00*S3+(-5.978055e+00)*S4+(-3.797963e+00)*S5+(-4.035935e+00)*S6+1.057841e+00*S7+(-1.490302e+01)*S8+(-1.850793e+00)*S9 \
V2_part2=V2_part1+9.739863e-01*S10+0.000000e+00*S11+(-1.196249e+01)*S12+1.871138e+00*S13+2.847095e+00*S14+2.187812e+00*S15+0.000000e+00*S16+4.250641e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V2_part3=V2_part2+(-1.111248e+00)*S20+0.000000e+00*S21+4.677533e+00*S22+0.000000e+00*S23+8.551933e+00*S24+1.180495e+01*S25+0.000000e+00*S26+0.000000e+00*S27+7.109069e-02*S28+3.542413e+00*S29 \
V2_part4=V2_part3+4.598689e+00*S30+1.688026e+01*S31+0.000000e+00*S32+1.608726e+00*S33+(-2.887320e+00)*S34+(-5.498282e-01)*S35+0.000000e+00*S36+0.000000e+00*S37+7.185200e+00*S38+1.200065e+00*S39 \
V2=V2_part4+0.000000e+00*S40+1.624581e-01*S41 \
V3_part1=(-5.086318e-01)*S0+(-1.666454e+00)*S1+6.551478e-01*S2+7.926928e-01*S3+(-9.036834e-01)*S4+(-6.401197e-01)*S5+(-9.219478e-01)*S6+2.141287e+00*S7+(-1.866846e+00)*S8+(-6.234483e-01)*S9 \
V3_part2=V3_part1+(-1.078128e-01)*S10+(-1.890887e+00)*S11+(-5.321143e+00)*S12+(-1.471397e+00)*S13+(-1.758897e+00)*S14+(-3.694665e-01)*S15+3.970089e-01*S16+(-1.033010e+00)*S17+(-1.301655e+00)*S18+(-2.864516e+00)*S19 \
V3_part3=V3_part2+(-5.853030e-01)*S20+(-1.470865e+00)*S21+(-2.616547e+00)*S22+(-9.327788e-01)*S23+(-2.212609e+00)*S24+(-2.543063e+00)*S25+(-5.770013e+00)*S26+(-4.621301e-01)*S27+(-1.014467e+00)*S28+6.510957e-01*S29 \
V3_part4=V3_part3+(-2.413413e+00)*S30+(-2.717566e+00)*S31+(-3.993186e+01)*S32+(-1.848928e-01)*S33+(-5.032748e+00)*S34+(-5.964708e+00)*S35+(-8.191784e-01)*S36+(-2.217119e+00)*S37+(-1.082177e+01)*S38+(-6.118943e-02)*S39 \
V3=V3_part4+(-1.198752e+00)*S40+(-5.100407e+01)*S41 \
V4_part1=(-3.030746e-01)*S0+4.757088e+00*S1+(-1.036001e+00)*S2+(-2.008637e+00)*S3+1.897272e+00*S4+3.190063e+00*S5+1.017682e+00*S6+(-3.648642e+00)*S7+2.981893e+00*S8+1.133451e+00*S9 \
V4_part2=V4_part1+(-1.062747e+00)*S10+(-9.976251e-01)*S11+9.128155e+00*S12+7.644196e+00*S13+4.710130e+00*S14+1.587099e+00*S15+(-1.018012e+00)*S16+2.113388e+00*S17+8.822365e+00*S18+8.928717e+00*S19 \
V4_part3=V4_part2+2.841530e-02*S20+9.000384e+00*S21+8.280415e+00*S22+4.526142e-02*S23+1.672246e+01*S24+1.008850e+01*S25+1.136563e+01*S26+(-9.185324e-01)*S27+(-5.170789e-01)*S28+(-2.522778e+00)*S29 \
V4_part4=V4_part3+2.014585e+01*S30+1.146195e+01*S31+8.469307e+01*S32+1.071761e+00*S33+1.808034e+01*S34+1.155876e+01*S35+1.460057e+01*S36+1.207637e+01*S37+2.156946e+01*S38+1.421376e+00*S39 \
V4=V4_part4+4.281367e+00*S40+1.079896e+02*S41 \
V5_part1=2.003511e+00*S0+5.398670e-01*S1+5.278480e+00*S2+3.722306e+00*S3+7.065587e-01*S4+2.406223e-01*S5+1.102692e+00*S6+1.017270e+01*S7+5.828565e-01*S8+5.616177e-01*S9 \
V5_part2=V5_part1+2.042986e+00*S10+3.843229e+00*S11+1.147986e+00*S12+4.282797e-01*S13+6.276933e-01*S14+4.952102e-01*S15+2.390050e+00*S16+8.181928e-01*S17+5.413850e-01*S18+9.059899e-01*S19 \
V5_part3=V5_part2+3.193236e+00*S20+4.876243e-01*S21+7.530507e-01*S22+2.956425e+00*S23+7.212123e-01*S24+9.848546e-01*S25+1.637893e+00*S26+3.017612e+00*S27+3.712150e+00*S28+4.748411e+00*S29 \
V5_part4=V5_part3+8.641450e-01*S30+1.185907e+00*S31+1.876870e+00*S32+2.499326e+00*S33+1.170749e+00*S34+1.713536e+00*S35+8.088107e-01*S36+1.279248e+00*S37+2.646765e+00*S38+3.006074e+00*S39 \
V5=V5_part4+1.479734e+00*S40+1.771278e+00*S41 \
V6_part1=5.631525e-02*S0+(-4.527483e-02)*S1+2.433467e-01*S2+1.988157e-01*S3+(-8.611867e-02)*S4+(-1.012093e-02)*S5+(-3.492312e-03)*S6+7.762928e-03*S7+(-5.495205e-02)*S8+(-6.935987e-02)*S9 \
V6_part2=V6_part1+6.653515e-02*S10+1.177488e-01*S11+(-2.575131e-01)*S12+(-3.753328e-02)*S13+(-4.941885e-02)*S14+(-5.138858e-02)*S15+1.770887e-01*S16+(-1.111095e-01)*S17+(-4.744182e-02)*S18+(-1.208638e-01)*S19 \
V6_part3=V6_part2+1.814210e-01*S20+(-5.566582e-02)*S21+(-1.316751e-01)*S22+2.369172e-01*S23+(-1.108639e-01)*S24+(-1.685893e-01)*S25+(-3.214993e-01)*S26+8.615794e-02*S27+1.460738e-01*S28+2.063744e-01*S29 \
V6_part4=V6_part3+(-1.107837e-01)*S30+(-1.865126e-01)*S31+(-1.331928e+00)*S32+8.865362e-02*S33+(-2.920246e-01)*S34+(-3.646315e-01)*S35+(-5.748482e-02)*S36+(-2.295430e-01)*S37+(-6.769526e-01)*S38+1.652510e-01*S39 \
V6=V6_part4+1.350984e-01*S40+(-1.670347e+00)*S41 \
V7_part1=1.177837e+00*S0+1.500517e+00*S1+1.206774e+00*S2+1.396366e+00*S3+1.503262e+00*S4+7.683736e-01*S5+8.130756e-01*S6+1.299806e+00*S7+9.784926e-01*S8+9.152801e-01*S9 \
V7_part2=V7_part1+2.163132e+00*S10+2.420000e+00*S11+3.128094e+00*S12+1.801319e+00*S13+1.931912e+00*S14+1.692363e+00*S15+1.745893e+00*S16+1.900407e+00*S17+3.822121e+00*S18+4.258233e+00*S19 \
V7_part3=V7_part2+4.090153e+00*S20+2.960161e+00*S21+3.302354e+00*S22+3.145160e+00*S23+5.642279e+00*S24+6.021139e+00*S25+6.552591e+00*S26+3.919923e+00*S27+4.360751e+00*S28+4.634215e+00*S29 \
V7_part4=V7_part3+7.508414e+00*S30+8.023023e+00*S31+1.050508e+01*S32+5.551362e+00*S33+6.992797e+00*S34+7.348933e+00*S35+9.519923e+00*S36+1.034105e+01*S37+1.156421e+01*S38+7.410988e+00*S39 \
V7=V7_part4+8.248991e+00*S40+1.189972e+01*S41 \
V8_part1=(-4.715267e-02)*S0+1.982683e-02*S1+(-6.975446e-02)*S2+(-3.886189e-01)*S3+3.556227e-02*S4+(-2.627607e-02)*S5+(-9.510023e-02)*S6+1.881319e-02*S7+(-1.152053e-01)*S8+(-1.652407e-02)*S9 \
V8_part2=V8_part1+(-2.334803e-02)*S10+(-3.519434e-01)*S11+(-1.721717e-01)*S12+1.018985e-01*S13+(-4.721076e-02)*S14+9.118813e-02*S15+(-4.820438e-01)*S16+2.715558e-02*S17+5.262696e-01*S18+2.318731e-01*S19 \
V8_part3=V8_part2+(-9.310698e-01)*S20+2.982757e-01*S21+6.836660e-02*S22+(-9.768660e-01)*S23+1.175408e+00*S24+4.270604e-01*S25+(-2.767179e-01)*S26+1.137967e-01*S27+(-4.126207e-01)*S28+(-1.016600e+00)*S29 \
V8_part4=V8_part3+1.897734e+00*S30+8.511666e-01*S31+1.446960e+00*S32+4.400144e-01*S33+9.004568e-01*S34+(-3.574909e-01)*S35+2.298670e+00*S36+1.635055e+00*S37+6.863992e-01*S38+8.264228e-01*S39 \
V8=V8_part4+4.014904e-01*S40+1.749984e+00*S41 \
V9_part1=(-1.717418e+00)*S0+(-2.017413e+00)*S1+(-5.905404e-01)*S2+(-4.063957e+00)*S3+(-9.510243e-01)*S4+(-4.038184e+00)*S5+(-3.287736e+00)*S6+(-4.523870e-01)*S7+1.540071e-01*S8+(-1.298732e+00)*S9 \
V9_part2=V9_part1+(-2.937191e+00)*S10+(-4.084889e+00)*S11+(-1.390861e+00)*S12+(-9.819029e-01)*S13+(-1.172294e+00)*S14+5.093348e+00*S15+(-8.495621e+00)*S16+(-4.884634e-01)*S17+(-1.907840e+00)*S18+(-1.760308e+00)*S19 \
V9_part3=V9_part2+(-1.796663e+01)*S20+(-1.146444e+00)*S21+(-2.150855e+00)*S22+(-1.481382e+01)*S23+(-4.595518e-01)*S24+(-2.673887e-01)*S25+(-3.381815e-01)*S26+(-3.005108e+00)*S27+(-7.010928e+00)*S28+(-1.403414e+01)*S29 \
V9_part4=V9_part3+5.786383e-01*S30+1.361688e+00*S31+(-4.672337e+00)*S32+(-4.517269e+00)*S33+(-2.145476e+00)*S34+1.319207e-01*S35+7.803240e+00*S36+(-6.020467e+00)*S37+(-2.196372e+00)*S38+(-4.628485e+00)*S39 \
V9=V9_part4+1.896747e+03*S40+(-4.422523e+00)*S41 \
V10_part1=8.694189e+00*S0+1.054768e+00*S1+2.539367e+00*S2+6.430218e+00*S3+(-7.231204e-02)*S4+2.121441e+00*S5+9.049649e+00*S6+1.497272e+00*S7+(-3.678985e+00)*S8+7.425204e-01*S9 \
V10_part2=V10_part1+1.627143e+01*S10+1.270084e+01*S11+(-1.049018e+00)*S12+2.669643e+00*S13+(-1.003506e-01)*S14+(-1.275543e+01)*S15+1.389369e+01*S16+(-3.236992e-01)*S17+(-1.866835e+00)*S18+(-3.451867e+00)*S19 \
V10_part3=V10_part2+3.035694e+01*S20+(-7.256854e-01)*S21+(-1.713608e+00)*S22+2.473070e+01*S23+2.080585e+00*S24+(-9.190723e+00)*S25+(-5.324384e+00)*S26+2.141080e+01*S27+2.276356e+01*S28+2.417187e+01*S29 \
V10_part4=V10_part3+9.945069e-01*S30+(-1.447105e+01)*S31+6.948329e+00*S32+3.505252e+01*S33+8.888173e-01*S34+(-7.889358e+00)*S35+(-2.700995e+01)*S36+(-1.125594e+01)*S37+7.986244e-01*S38+4.138775e+01*S39 \
V10=V10_part4+1.000000e+04*S40+6.942141e+00*S41 \
V11_part1=6.725952e-01*S0+4.125275e+00*S1+9.403433e-01*S2+1.588626e+00*S3+7.328362e+00*S4+4.159952e+00*S5+9.656041e-01*S6+7.295611e-01*S7+5.656524e+00*S8+6.587562e+00*S9 \
V11_part2=V11_part1+9.319743e-01*S10+1.341250e+00*S11+6.291160e+00*S12+2.354042e+00*S13+5.079142e+00*S14+1.524896e+01*S15+1.991688e+00*S16+8.548745e+00*S17+6.830933e+00*S18+8.424714e+00*S19 \
V11_part3=V11_part2+3.399750e+00*S20+4.465901e+00*S21+6.553591e+00*S22+2.734796e+00*S23+4.656967e+00*S24+1.161692e+01*S25+1.255108e+01*S26+1.162807e+00*S27+1.943000e+00*S28+3.135614e+00*S29 \
V11_part4=V11_part3+5.516210e+00*S30+1.502682e+01*S31+5.243199e+00*S32+1.517829e+00*S33+7.052445e+00*S34+1.467726e+01*S35+1.195584e+01*S36+1.952713e+01*S37+1.179339e+01*S38+1.761307e+00*S39 \
V11=V11_part4+(-1.248414e+03)*S40+5.309289e+00*S41 \
V12_part1=(-2.660932e-02)*S0+8.198896e-02*S1+(-6.908388e-02)*S2+(-1.885490e-01)*S3+3.447068e-01*S4+3.892634e-01*S5+(-8.996558e-02)*S6+(-6.177082e-02)*S7+1.880000e-01*S8+1.335367e-01*S9 \
V12_part2=V12_part1+(-9.684939e-02)*S10+(-1.993905e-01)*S11+1.530545e-01*S12+(-1.076647e-02)*S13+1.652676e-01*S14+1.222985e+00*S15+(-1.974633e-01)*S16+4.405405e-01*S17+2.336561e-01*S18+4.862099e-01*S19 \
V12_part3=V12_part2+(-8.757832e-01)*S20+1.044843e-01*S21+1.253615e-01*S22+(-4.259687e-01)*S23+1.998825e-01*S24+(-1.911664e-02)*S25+(-5.579650e-01)*S26+(-1.490846e-01)*S27+(-3.797705e-01)*S28+(-6.268321e-01)*S29 \
V12_part4=V12_part3+3.925336e-01*S30+(-5.489720e-01)*S31+(-2.018091e-01)*S32+(-2.318114e-01)*S33+5.570398e-01*S34+(-6.435148e-01)*S35+(-3.196445e-01)*S36+(-7.797165e-01)*S37+(-5.737704e-01)*S38+(-2.515311e-01)*S39 \
V12=V12_part4+2.075174e+00*S40+(-4.815890e-02)*S41 \
V13_part1=2.667890e+00*S0+2.628690e+00*S1+2.661218e+00*S2+3.320718e+00*S3+2.479056e+00*S4+1.236309e+00*S5+1.905595e+00*S6+1.595152e+00*S7+1.600104e+00*S8+1.661757e+00*S9 \
V13_part2=V13_part1+5.020778e+00*S10+5.521585e+00*S11+5.246023e+00*S12+3.159285e+00*S13+3.408502e+00*S14+2.472141e+00*S15+4.273476e+00*S16+3.170123e+00*S17+6.780892e+00*S18+7.417044e+00*S19 \
V13_part3=V13_part2+9.981425e+00*S20+5.207884e+00*S21+5.697314e+00*S22+7.557322e+00*S23+9.840692e+00*S24+1.056979e+01*S25+1.192782e+01*S26+8.838797e+00*S27+9.946925e+00*S28+1.078287e+01*S29 \
V13_part4=V13_part3+1.312917e+01*S30+1.468746e+01*S31+1.633163e+01*S32+1.257148e+01*S33+1.199184e+01*S34+1.359381e+01*S35+1.719805e+01*S36+1.868559e+01*S37+2.075702e+01*S38+1.651392e+01*S39 \
V13=V13_part4+1.165652e+01*S40+1.793006e+01*S41 \
V14_part1=1.792446e-01*S0+(-2.797906e-01)*S1+1.721547e-01*S2+(-3.132773e-01)*S3+(-3.037243e-01)*S4+(-2.790292e-01)*S5+(-3.639027e-02)*S6+2.113766e-02*S7+(-4.538105e-01)*S8+(-2.150934e-01)*S9 \
V14_part2=V14_part1+5.409948e-01*S10+1.041204e-01*S11+(-1.239043e+00)*S12+(-6.050136e-02)*S13+(-5.145312e-01)*S14+(-5.156739e-01)*S15+(-3.644340e-01)*S16+(-4.250734e-01)*S17+1.199534e-01*S18+(-9.813550e-01)*S19 \
V14_part3=V14_part2+(-7.440244e-02)*S20+(-7.488139e-02)*S21+(-5.811711e-01)*S22+(-5.227632e-01)*S23+7.747861e-01*S24+6.176280e-02*S25+(-1.305903e+00)*S26+1.287240e+00*S27+6.805945e-01*S28+(-5.608583e-01)*S29 \
V14_part4=V14_part3+1.547436e+00*S30+8.415287e-01*S31+(-1.298275e+00)*S32+2.569185e+00*S33+(-7.736323e-01)*S34+(-1.858228e+00)*S35+3.400983e+00*S36+2.273860e+00*S37+(-9.743534e-01)*S38+4.116880e+00*S39 \
V14=V14_part4+3.591168e+00*S40+(-1.554375e+00)*S41 \
V15_part1=(-6.987656e-02)*S0+1.246145e-01*S1+1.497354e-02*S2+3.197761e-01*S3+(-8.121122e-03)*S4+(-2.309045e-01)*S5+9.810540e-01*S6+1.249692e-01*S7+(-6.676595e-01)*S8+4.804826e-01*S9 \
V15_part2=V15_part1+(-1.590232e-02)*S10+(-1.553526e-02)*S11+(-2.874190e-01)*S12+5.383757e-01*S13+(-2.529597e-02)*S14+(-4.491553e-01)*S15+(-5.923750e-01)*S16+(-6.665634e-02)*S17+(-1.007932e-01)*S18+(-4.201404e-01)*S19 \
V15_part3=V15_part2+3.061282e-02*S20+(-2.041420e-01)*S21+(-4.660615e-01)*S22+(-4.069138e-01)*S23+1.229879e-01*S24+(-2.794097e+00)*S25+1.000000e+04*S26+(-5.501221e-02)*S27+(-2.883123e-01)*S28+(-1.994681e+00)*S29 \
V15_part4=V15_part3+(-1.021942e-01)*S30+7.028479e+00*S31+(-3.127637e-01)*S32+(-5.564608e-03)*S33+(-9.103866e-01)*S34+1.544111e+00*S35+8.439489e+03*S36+1.762965e+02*S37+3.687834e+03*S38+(-9.304354e-02)*S39 \
V15=V15_part4+2.779389e+00*S40+(-4.190920e-01)*S41 \
V16_part1=3.309467e+00*S0+2.919271e+00*S1+6.203802e-01*S2+7.344895e-01*S3+9.416089e-01*S4+3.136172e+00*S5+1.587015e+00*S6+9.774167e-02*S7+2.371347e+00*S8+2.684916e-01*S9 \
V16_part2=V16_part1+4.050896e+00*S10+2.323685e+00*S11+2.728838e+00*S12+3.015499e+00*S13+1.668837e+00*S14+1.151923e+00*S15+2.106691e+00*S16+1.013106e+00*S17+4.226440e+00*S18+3.027336e+00*S19 \
V16_part3=V16_part2+1.907629e+00*S20+5.749119e+00*S21+4.355630e+00*S22+1.619885e+00*S23+5.033858e+00*S24+1.251476e+01*S25+1.000000e+04*S26+5.450383e+00*S27+3.058713e+00*S28+5.176178e+00*S29 \
V16_part4=V16_part3+5.935325e+00*S30+6.988521e+03*S31+3.226272e+00*S32+5.962892e+00*S33+4.247930e+00*S34+2.667994e+02*S35+1.000000e+04*S36+5.318094e+03*S37+5.411062e+03*S38+5.933919e+00*S39 \
V16=V16_part4+(-1.121310e-01)*S40+2.826829e+00*S41 \
V17_part1=1.977424e-02*S0+(-4.463844e-01)*S1+(-1.872871e-02)*S2+(-1.926739e-01)*S3+8.381555e-02*S4+7.854339e-01*S5+(-2.961904e-01)*S6+(-2.295837e-01)*S7+2.534870e-01*S8+(-1.421364e-01)*S9 \
V17_part2=V17_part1+6.596971e-02*S10+4.625138e-01*S11+1.629313e-01*S12+1.457026e-01*S13+2.684311e-01*S14+1.491675e-01*S15+2.800601e-01*S16+6.478704e-02*S17+3.478841e-01*S18+8.396566e-01*S19 \
V17_part3=V17_part2+5.688145e-01*S20+1.249388e-01*S21+5.569618e-01*S22+7.257082e-01*S23+6.015313e-01*S24+3.395775e+00*S25+1.000000e+04*S26+(-6.208479e-02)*S27+1.032885e+00*S28+9.478172e-01*S29 \
V17_part4=V17_part3+8.315672e-01*S30+4.016693e+01*S31+1.843211e+00*S32+5.226954e-01*S33+1.965469e+00*S34+4.674854e+00*S35+9.778232e+03*S36+8.270737e+01*S37+9.512410e+03*S38+1.198781e+00*S39 \
V17=V17_part4+(-7.226616e+00)*S40+2.501541e+00*S41 \
V18_part1=(-5.887770e-01)*S0+1.372473e-01*S1+(-1.843420e+00)*S2+(-1.537212e+00)*S3+(-5.424415e-01)*S4+(-1.770101e+00)*S5+(-2.280052e-01)*S6+(-1.756822e+00)*S7+(-1.424440e-02)*S8+1.636170e-01*S9 \
V18_part2=V18_part1+(-4.917644e-01)*S10+(-1.100149e+00)*S11+7.493194e-02*S12+(-4.151920e-01)*S13+(-1.892340e+00)*S14+(-1.020647e+00)*S15+(-1.636209e+00)*S16+(-6.841548e-01)*S17+(-4.468054e-01)*S18+(-1.353818e+00)*S19 \
V18_part3=V18_part2+(-8.270951e-01)*S20+(-3.215343e-01)*S21+(-1.561817e-01)*S22+(-2.007888e+00)*S23+1.697946e-01*S24+(-3.823415e-01)*S25+(-1.613210e+00)*S26+(-4.726178e-01)*S27+(-7.994281e-01)*S28+(-1.187359e+00)*S29 \
V18_part4=V18_part3+1.362573e-01*S30+(-1.146605e+00)*S31+(-9.839759e-01)*S32+(-9.678536e-02)*S33+(-7.137705e-01)*S34+(-1.248213e+00)*S35+(-6.878179e-01)*S36+(-1.761714e+00)*S37+(-1.428053e+00)*S38+(-2.823769e-01)*S39 \
V18=V18_part4+(-1.159097e+00)*S40+5.010843e-01*S41 \
V19_part1=4.146024e+00*S0+5.924397e-01*S1+5.171319e+00*S2+4.481811e+00*S3+1.094357e+00*S4+8.896627e+00*S5+8.591735e-01*S6+5.506999e+00*S7+5.428364e-01*S8+6.232786e-01*S9 \
V19_part2=V19_part1+4.428165e+00*S10+5.444593e+00*S11+1.199455e+00*S12+4.143428e+00*S13+5.554711e+00*S14+2.088280e+00*S15+5.524961e+00*S16+9.368550e-01*S17+4.680333e+00*S18+5.688731e+00*S19 \
V19_part3=V19_part2+3.070352e+00*S20+4.944452e+00*S21+1.872321e+00*S22+5.584036e+00*S23+4.966507e-01*S24+1.944913e+00*S25+6.082092e+00*S26+4.833544e+00*S27+3.286908e+00*S28+4.387951e+00*S29 \
V19_part4=V19_part3+1.287282e+00*S30+6.259055e+00*S31+5.162123e+00*S32+1.623817e+00*S33+2.532314e+00*S34+3.226537e+00*S35+6.943132e+00*S36+8.074998e+00*S37+3.445796e+00*S38+2.266470e+00*S39 \
V19=V19_part4+6.143244e+00*S40+2.868959e+00*S41 \
V20_part1=3.747349e+00*S0+3.118365e+00*S1+5.728398e+00*S2+5.718643e+00*S3+7.333462e+00*S4+5.158837e+00*S5+3.039084e+00*S6+3.557307e+00*S7+5.263491e+00*S8+5.018063e+00*S9 \
V20_part2=V20_part1+5.019531e+00*S10+6.346003e+00*S11+8.087696e+00*S12+3.815832e+00*S13+5.779771e+00*S14+5.802684e+00*S15+6.080722e+00*S16+5.316421e+00*S17+7.161827e+00*S18+8.529672e+00*S19 \
V20_part3=V20_part2+8.425571e+00*S20+5.305941e+00*S21+3.903387e+00*S22+9.228752e+00*S23+5.848963e+00*S24+5.115106e+00*S25+7.358388e+00*S26+7.556930e+00*S27+7.202864e+00*S28+6.922260e+00*S29 \
V20_part4=V20_part3+8.466449e+00*S30+4.804728e+00*S31+1.053569e+01*S32+7.307389e+00*S33+8.857286e+00*S34+7.617362e+00*S35+9.653698e+00*S36+1.560539e+01*S37+1.037075e+01*S38+8.616758e+00*S39 \
V20=V20_part4+9.555857e+00*S40+1.083756e+01*S41 \
V21_part1=6.915189e+00*S0+7.331395e+00*S1+9.110092e+00*S2+4.492393e+00*S3+(-4.234110e+00)*S4+2.244568e+01*S5+4.095575e+00*S6+4.886069e+00*S7+6.078937e+00*S8+(-5.288506e+00)*S9 \
V21_part2=V21_part1+6.955392e+00*S10+9.937072e+00*S11+5.230892e+00*S12+1.502986e+01*S13+(-2.349116e+01)*S14+6.825789e+00*S15+2.968042e+03*S16+6.406017e+00*S17+6.014438e+00*S18+8.187932e+00*S19 \
V21_part3=V21_part2+2.369511e+00*S20+1.249079e+01*S21+2.198440e+00*S22+5.525758e+00*S23+1.030683e+01*S24+0.000000e+00*S25+2.181737e+00*S26+6.277607e+00*S27+2.589256e+00*S28+(-9.792126e+01)*S29 \
V21_part4=V21_part3+6.322859e+00*S30+2.636722e+00*S31+2.414287e+00*S32+6.722077e+00*S33+7.329921e+00*S34+3.415813e+01*S35+(-1.988893e+03)*S36+(-2.404849e+02)*S37+0.000000e+00*S38+8.669432e+00*S39 \
V21=V21_part4+2.558385e+00*S40+1.571993e+00*S41 \
V22_part1=(-3.483333e+00)*S0+1.898328e+00*S1+(-1.312035e+00)*S2+(-1.384794e+00)*S3+7.314464e+00*S4+(-2.547182e+00)*S5+(-2.241936e+00)*S6+(-1.442399e+00)*S7+(-2.970398e+00)*S8+1.152042e+01*S9 \
V22_part2=V22_part1+(-3.678434e+00)*S10+(-3.779810e+00)*S11+(-2.217342e+00)*S12+(-2.104052e+00)*S13+3.025339e+01*S14+(-2.642014e+00)*S15+8.859840e+03*S16+(-1.963032e+00)*S17+(-5.160090e+00)*S18+2.922120e-01*S19 \
V22_part3=V22_part2+(-1.117392e+00)*S20+(-1.307845e+01)*S21+(-1.852110e+00)*S22+(-6.255228e-02)*S23+(-8.882255e-01)*S24+0.000000e+00*S25+(-1.062622e+00)*S26+(-6.628970e+00)*S27+(-7.875882e-01)*S28+5.656420e+00*S29 \
V22_part4=V22_part3+(-1.559899e+00)*S30+(-1.249561e+00)*S31+(-1.426571e+00)*S32+(-1.679098e+00)*S33+(-1.794376e+00)*S34+9.246203e-01*S35+5.867440e-01*S36+(-1.555047e+01)*S37+0.000000e+00*S38+(-8.044205e-01)*S39 \
V22=V22_part4+(-1.556490e+00)*S40+(-9.646265e-01)*S41 \
V23_part1=(-4.336605e+00)*S0+(-7.774619e+00)*S1+(-4.806445e+00)*S2+(-1.837791e+00)*S3+5.768229e+00*S4+(-1.694428e+01)*S5+(-1.651647e+00)*S6+(-1.790837e+00)*S7+(-2.748443e+00)*S8+4.231575e+00*S9 \
V23_part2=V23_part1+(-6.212400e+00)*S10+(-9.460647e+00)*S11+(-3.238888e+00)*S12+(-1.312741e+01)*S13+5.813071e+01*S14+(-2.518710e+00)*S15+(-1.000000e+04)*S16+(-1.549532e+00)*S17+(-3.823614e+00)*S18+(-9.965619e+00)*S19 \
V23_part3=V23_part2+3.611024e-01*S20+(-7.639561e+00)*S21+1.821928e+00*S22+(-6.197374e+00)*S23+(-1.303649e+01)*S24+0.000000e+00*S25+(-4.888095e-01)*S26+(-2.904555e+00)*S27+9.255488e-01*S28+4.951690e+02*S29 \
V23_part4=V23_part3+(-6.240775e+00)*S30+(-2.093814e+00)*S31+7.408199e-01*S32+(-6.925575e+00)*S33+(-7.662316e+00)*S34+(-6.514999e+01)*S35+1.000000e+04*S36+1.426854e+03*S37+0.000000e+00*S38+(-1.217017e+01)*S39 \
V23=V23_part4+6.816665e-01*S40+2.292312e+01*S41 \
V24_part1=6.770968e+00*S0+1.034119e+01*S1+0.000000e+00*S2+1.613178e+01*S3+7.894874e+01*S4+(-2.704753e+00)*S5+0.000000e+00*S6+1.278212e+01*S7+3.314696e+01*S8+7.514605e+01*S9 \
V24_part2=V24_part1+4.796571e+00*S10+3.425297e+01*S11+(-1.468045e+01)*S12+1.877269e+01*S13+2.325898e+01*S14+8.959182e+00*S15+(-7.216639e+00)*S16+1.325118e+01*S17+1.263457e+01*S18+0.000000e+00*S19 \
V24_part3=V24_part2+2.726242e+01*S20+2.390064e+00*S21+2.207319e+01*S22+(-3.141448e+01)*S23+2.281008e+00*S24+3.958468e+02*S25+1.039196e+01*S26+4.448053e+00*S27+2.784208e+01*S28+4.494289e+01*S29 \
V24_part4=V24_part3+1.197937e+01*S30+(-2.511617e+02)*S31+(-1.828402e+01)*S32+2.283975e+00*S33+(-1.319434e+01)*S34+(-1.907199e+02)*S35+4.827614e+00*S36+(-2.003825e+01)*S37+0.000000e+00*S38+(-2.157970e+01)*S39 \
V24=V24_part4+(-2.049606e+00)*S40+(-1.090408e+02)*S41 \
V25_part1=6.209722e+01*S0+1.710260e+01*S1+0.000000e+00*S2+5.797455e+01*S3+(-5.425656e+01)*S4+3.587205e+01*S5+0.000000e+00*S6+4.264043e+01*S7+1.793355e+01*S8+(-6.142632e+01)*S9 \
V25_part2=V25_part1+8.256113e+01*S10+4.253037e+01*S11+2.386011e+01*S12+7.205535e+01*S13+4.815801e+01*S14+3.282120e+01*S15+9.046279e+01*S16+1.561034e+01*S17+1.186976e+02*S18+0.000000e+00*S19 \
V25_part3=V25_part2+9.847829e+01*S20+1.106334e+02*S21+4.311109e+01*S22+(-4.369783e+00)*S23+6.167934e+01*S24+1.554355e+02*S25+8.157809e+01*S26+1.322613e+02*S27+5.346422e+01*S28+3.794378e+01*S29 \
V25_part4=V25_part3+7.888713e+01*S30+2.192205e+02*S31+4.998983e+01*S32+1.062231e+02*S33+1.137464e+02*S34+1.716115e+02*S35+8.386562e+01*S36+8.121020e+01*S37+0.000000e+00*S38+1.521192e+02*S39 \
V25=V25_part4+9.655525e+01*S40+1.804284e+02*S41 \
V26_part1=2.417700e+01*S0+2.385171e+01*S1+0.000000e+00*S2+1.134307e+00*S3+1.733718e+01*S4+2.205910e+01*S5+0.000000e+00*S6+1.885839e+01*S7+1.237649e+01*S8+1.842793e+01*S9 \
V26_part2=V26_part1+3.575944e+01*S10+4.668927e+00*S11+3.860090e+01*S12+1.371709e+01*S13+1.036178e+01*S14+2.569648e+01*S15+2.108200e+01*S16+2.456511e+01*S17+1.800807e+01*S18+0.000000e+00*S19 \
V26_part3=V26_part2+6.409454e+00*S20+3.957173e+01*S21+(-2.045836e+01)*S22+2.071010e+02*S23+3.763846e+01*S24+(-2.857685e+02)*S25+1.889456e+02*S26+2.161054e+01*S27+4.985611e+00*S28+1.219230e+02*S29 \
V26_part4=V26_part3+3.625185e+01*S30+1.258563e+03*S31+2.924938e+02*S32+3.618645e+01*S33+3.571393e+01*S34+1.060985e+03*S35+1.776725e+02*S36+9.927335e+01*S37+0.000000e+00*S38+1.454710e+02*S39 \
V26=V26_part4+1.722056e+02*S40+3.247916e+02*S41 \
V27_part1=(-5.669178e-01)*S0+(-1.172038e-01)*S1+(-1.953953e+00)*S2+(-1.836642e+00)*S3+(-5.620303e-01)*S4+(-1.633308e+00)*S5+(-3.993366e-01)*S6+(-1.998826e+00)*S7+(-4.672230e-01)*S8+1.326299e-01*S9 \
V27_part2=V27_part1+(-5.094759e-01)*S10+(-1.433521e+00)*S11+(-8.730346e-02)*S12+(-5.554674e-01)*S13+(-2.113030e+00)*S14+(-1.299838e+00)*S15+(-1.892630e+00)*S16+(-8.769771e-01)*S17+(-7.448242e-01)*S18+(-1.651374e+00)*S19 \
V27_part3=V27_part2+(-1.009859e+00)*S20+(-3.133706e-01)*S21+(-2.833434e-01)*S22+(-2.085954e+00)*S23+4.230250e-02*S24+(-5.268507e-01)*S25+(-1.734025e+00)*S26+(-8.274065e-01)*S27+(-1.045979e+00)*S28+(-1.424241e+00)*S29 \
V27_part4=V27_part3+(-1.445632e-01)*S30+(-1.389897e+00)*S31+(-1.026876e+00)*S32+(-2.895915e-01)*S33+(-9.836223e-01)*S34+(-1.792708e+00)*S35+(-4.728656e-01)*S36+(-1.421940e+00)*S37+(-1.789996e+00)*S38+(-5.703434e-01)*S39 \
V27=V27_part4+(-1.507365e+00)*S40+3.616808e-01*S41 \
V28_part1=4.115322e+00*S0+1.274062e+00*S1+5.077989e+00*S2+4.593521e+00*S3+9.607968e-01*S4+8.096580e+00*S5+6.888639e-01*S6+5.873685e+00*S7+9.056959e-01*S8+5.504149e-01*S9 \
V28_part2=V28_part1+4.146317e+00*S10+5.527164e+00*S11+1.389632e+00*S12+3.913677e+00*S13+5.651624e+00*S14+2.046285e+00*S15+5.633764e+00*S16+1.046053e+00*S17+4.733265e+00*S18+5.844260e+00*S19 \
V28_part3=V28_part2+3.037742e+00*S20+4.984088e+00*S21+1.814966e+00*S22+5.301949e+00*S23+4.862436e-02*S24+2.056178e+00*S25+6.096137e+00*S26+6.141480e+00*S27+3.346519e+00*S28+4.628941e+00*S29 \
V28_part4=V28_part3+1.108043e+00*S30+6.190611e+00*S31+5.080918e+00*S32+1.204686e+00*S33+2.331390e+00*S34+3.561676e+00*S35+5.804731e+00*S36+6.561947e+00*S37+3.676765e+00*S38+1.527308e+00*S39 \
V28=V28_part4+5.898771e+00*S40+2.859922e+00*S41 \
V29_part1=3.745485e+00*S0+3.121798e+00*S1+6.005981e+00*S2+6.506750e+00*S3+7.580853e+00*S4+4.932745e+00*S5+3.625157e+00*S6+3.754990e+00*S7+5.539637e+00*S8+5.264200e+00*S9 \
V29_part2=V29_part1+5.025924e+00*S10+6.889892e+00*S11+7.561165e+00*S12+4.064928e+00*S13+6.059702e+00*S14+6.139521e+00*S15+6.236867e+00*S16+5.420825e+00*S17+7.217682e+00*S18+8.060001e+00*S19 \
V29_part3=V29_part2+8.146377e+00*S20+4.417655e+00*S21+3.813872e+00*S22+9.314925e+00*S23+5.672221e+00*S24+4.152497e+00*S25+6.250906e+00*S26+6.688829e+00*S27+6.939233e+00*S28+6.007922e+00*S29 \
V29_part4=V29_part3+8.224598e+00*S30+4.189454e+00*S31+9.452493e+00*S32+7.008911e+00*S33+8.583242e+00*S34+6.610723e+00*S35+6.656870e+00*S36+8.368112e+00*S37+8.603434e+00*S38+8.417987e+00*S39 \
V29=V29_part4+9.745466e+00*S40+9.594347e+00*S41 \
V30_part1=4.266101e-01*S0+6.028985e+00*S1+7.053132e+00*S2+7.581430e+00*S3+(-9.916929e+00)*S4+2.215142e+02*S5+(-1.012971e+00)*S6+6.212836e+00*S7+2.085933e+01*S8+1.079765e+01*S9 \
V30_part2=V30_part1+1.296696e+01*S10+1.131879e+02*S11+6.692282e+00*S12+1.600348e+01*S13+6.399932e+00*S14+4.550194e+01*S15+9.513484e+00*S16+3.428197e+01*S17+1.000000e+04*S18+1.174020e+01*S19 \
V30_part3=V30_part2+1.315954e+01*S20+8.971787e+01*S21+2.197366e+01*S22+9.891905e+00*S23+(-3.713527e+01)*S24+5.360450e+02*S25+1.000000e+04*S26+1.857427e+01*S27+8.332477e+02*S28+5.978280e+03*S29 \
V30_part4=V30_part3+7.820882e+03*S30+1.341267e+03*S31+(-3.831761e+01)*S32+8.662248e+00*S33+(-4.674742e+02)*S34+4.455233e-01*S35+(-1.716639e+03)*S36+(-1.943263e+02)*S37+1.999128e+01*S38+5.682364e+00*S39 \
V30=V30_part4+2.463930e+01*S40+3.030808e+01*S41 \
V31_part1=2.103631e+02*S0+(-1.767406e+00)*S1+(-4.035268e+00)*S2+(-1.962669e+00)*S3+3.690290e+00*S4+3.611054e+01*S5+(-6.884313e+00)*S6+(-2.188861e+00)*S7+(-1.175961e+01)*S8+1.193255e+00*S9 \
V31_part2=V31_part1+(-1.267477e+01)*S10+2.169197e+01*S11+(-4.627635e+00)*S12+(-2.089012e+01)*S13+(-1.843134e+00)*S14+(-1.733396e+01)*S15+(-3.598765e+00)*S16+(-7.144884e+00)*S17+(-2.886452e+03)*S18+(-8.835750e+00)*S19 \
V31_part3=V31_part2+(-8.564134e+00)*S20+(-1.036134e+02)*S21+(-9.227445e+00)*S22+(-5.628872e+00)*S23+1.381957e+02*S24+(-6.854905e+01)*S25+1.000000e+04*S26+(-1.835596e+00)*S27+(-4.614273e+02)*S28+(-5.239650e+03)*S29 \
V31_part4=V31_part3+(-1.000000e+04)*S30+(-1.549104e+02)*S31+(-1.227208e+02)*S32+(-9.860275e+00)*S33+2.813221e+02*S34+2.465653e+00*S35+(-1.923511e+02)*S36+(-2.569518e+01)*S37+1.134016e+01*S38+(-6.325345e+00)*S39 \
V31=V31_part4+(-1.991668e+01)*S40+(-3.644762e+01)*S41 \
V32_part1=1.173481e+02*S0+(-4.190818e+00)*S1+(-1.554096e+00)*S2+(-4.419018e+00)*S3+3.095006e+01*S4+(-1.879002e+02)*S5+3.979180e+01*S6+(-1.940670e+00)*S7+(-3.757832e+00)*S8+(-6.611380e+00)*S9 \
V32_part2=V32_part1+(-4.947702e+00)*S10+(-1.832476e+02)*S11+1.460942e+01*S12+(-1.645735e+00)*S13+(-3.126210e+00)*S14+(-2.459949e+01)*S15+(-5.355508e+00)*S16+(-2.234325e+01)*S17+(-3.783429e+03)*S18+(-3.738077e+00)*S19 \
V32_part3=V32_part2+1.321184e+00*S20+2.372194e+02*S21+(-2.284145e+01)*S22+(-1.969002e+00)*S23+1.908004e+02*S24+(-1.030453e+02)*S25+1.000000e+04*S26+(-2.557406e+01)*S27+1.000000e+04*S28+1.741262e+03*S29 \
V32_part4=V32_part3+1.842546e+02*S30+(-2.220323e+03)*S31+1.932254e+03*S32+(-2.352087e+00)*S33+1.841059e+03*S34+1.062898e+03*S35+1.000000e+04*S36+1.150236e+03*S37+(-4.930587e+01)*S38+(-1.989003e+00)*S39 \
V32=V32_part4+(-8.818165e+00)*S40+1.196656e+02*S41 \
V33_part1=1.897607e+01*S0+0.000000e+00*S1+1.345056e+01*S2+0.000000e+00*S3+6.060170e+01*S4+(-3.201291e+00)*S5+1.368673e+01*S6+(-5.673480e-01)*S7+0.000000e+00*S8+6.115683e+01*S9 \
V33_part2=V33_part1+1.541053e+01*S10+(-2.036356e+01)*S11+0.000000e+00*S12+8.691001e+00*S13+1.200615e+01*S14+0.000000e+00*S15+(-4.514848e+00)*S16+0.000000e+00*S17+4.479953e+00*S18+0.000000e+00*S19 \
V33_part3=V33_part2+0.000000e+00*S20+1.373866e+01*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V33_part4=V33_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+6.353722e+00*S34+(-4.733055e+01)*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+4.256082e-01*S39 \
V33=V33_part4+0.000000e+00*S40+0.000000e+00*S41 \
V34_part1=1.012128e+01*S0+0.000000e+00*S1+2.511025e+01*S2+0.000000e+00*S3+(-5.528235e+01)*S4+3.824153e+01*S5+(-9.521448e+00)*S6+2.808082e+01*S7+0.000000e+00*S8+(-5.239096e+01)*S9 \
V34_part2=V34_part1+(-2.816060e+00)*S10+5.501967e+01*S11+0.000000e+00*S12+4.926842e-02*S13+2.551473e+01*S14+0.000000e+00*S15+4.210764e+01*S16+0.000000e+00*S17+(-1.773716e+01)*S18+0.000000e+00*S19 \
V34_part3=V34_part2+0.000000e+00*S20+(-2.045106e+01)*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V34_part4=V34_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+3.442046e+01*S34+1.414085e+02*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+5.549508e+01*S39 \
V34=V34_part4+0.000000e+00*S40+0.000000e+00*S41 \
V35_part1=(-3.154358e-01)*S0+0.000000e+00*S1+6.544827e+00*S2+0.000000e+00*S3+(-1.133626e+00)*S4+1.798052e+01*S5+7.217320e+00*S6+6.460546e+00*S7+0.000000e+00*S8+5.812401e+00*S9 \
V35_part2=V35_part1+6.665758e+00*S10+3.357616e+01*S11+0.000000e+00*S12+1.421786e+01*S13+6.644436e+00*S14+0.000000e+00*S15+8.817105e+00*S16+0.000000e+00*S17+2.960620e+01*S18+0.000000e+00*S19 \
V35_part3=V35_part2+0.000000e+00*S20+4.920773e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V35_part4=V35_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+5.946550e+01*S34+2.023991e+02*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+8.197461e+01*S39 \
V35=V35_part4+0.000000e+00*S40+0.000000e+00*S41 \
V36_part1=0.000000e+00*S0+(-2.461481e+00)*S1+0.000000e+00*S2+0.000000e+00*S3+(-6.054932e+00)*S4+0.000000e+00*S5+(-9.600224e-01)*S6+0.000000e+00*S7+(-2.860740e+00)*S8+(-5.219674e+00)*S9 \
V36_part2=V36_part1+0.000000e+00*S10+0.000000e+00*S11+(-4.018428e+00)*S12+0.000000e+00*S13+0.000000e+00*S14+(-2.248750e+00)*S15+0.000000e+00*S16+(-5.266116e+00)*S17+0.000000e+00*S18+0.000000e+00*S19 \
V36_part3=V36_part2+(-3.219135e+00)*S20+0.000000e+00*S21+(-2.562721e+00)*S22+0.000000e+00*S23+(-2.381533e+00)*S24+(-3.827788e+00)*S25+(-3.140539e+00)*S26+0.000000e+00*S27+(-2.435662e+00)*S28+(-3.260910e+00)*S29 \
V36_part4=V36_part3+(-3.086248e+00)*S30+(-3.703838e+00)*S31+(-6.142222e+00)*S32+(-2.361569e+00)*S33+(-3.086676e+00)*S34+(-3.212840e+00)*S35+(-3.730965e+00)*S36+(-4.646699e+00)*S37+(-6.889812e+00)*S38+(-2.669952e+00)*S39 \
V36=V36_part4+(-3.716073e+00)*S40+(-9.179857e+00)*S41 \
V37_part1=0.000000e+00*S0+8.266696e+00*S1+0.000000e+00*S2+0.000000e+00*S3+8.196344e+00*S4+0.000000e+00*S5+4.436906e+00*S6+0.000000e+00*S7+5.706020e+00*S8+7.518294e+00*S9 \
V37_part2=V37_part1+0.000000e+00*S10+0.000000e+00*S11+5.988314e+00*S12+0.000000e+00*S13+0.000000e+00*S14+6.129065e+00*S15+0.000000e+00*S16+8.029019e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V37_part3=V37_part2+4.224587e+00*S20+0.000000e+00*S21+5.081964e+00*S22+0.000000e+00*S23+9.427520e+00*S24+7.388505e+00*S25+1.190572e-01*S26+0.000000e+00*S27+4.688259e+00*S28+2.224768e+00*S29 \
V37_part4=V37_part3+9.483161e+00*S30+2.160727e+00*S31+3.504267e+00*S32+8.421607e+00*S33+7.348579e+00*S34+5.999018e+00*S35+1.381197e+00*S36+2.146783e+00*S37+8.893175e+00*S38+7.656733e+00*S39 \
V37=V37_part4+2.339835e+00*S40+8.458049e+00*S41 \
V38_part1=0.000000e+00*S0+2.025665e+00*S1+0.000000e+00*S2+0.000000e+00*S3+1.411698e+00*S4+0.000000e+00*S5+1.707748e+00*S6+0.000000e+00*S7+7.997423e-02*S8+8.756249e-01*S9 \
V38_part2=V38_part1+0.000000e+00*S10+0.000000e+00*S11+4.430749e+00*S12+0.000000e+00*S13+0.000000e+00*S14+2.265146e+00*S15+0.000000e+00*S16+7.413217e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V38_part3=V38_part2+8.431762e+00*S20+0.000000e+00*S21+9.661515e+00*S22+0.000000e+00*S23+8.877835e+00*S24+1.850881e+01*S25+1.844203e+01*S26+0.000000e+00*S27+8.383080e+00*S28+1.471613e+01*S29 \
V38_part4=V38_part3+9.605413e+00*S30+2.423932e+01*S31+2.021798e+01*S32+8.231038e+00*S33+1.068184e+01*S34+1.938396e+01*S35+2.006464e+01*S36+2.221695e+01*S37+2.917935e+01*S38+1.239730e+01*S39 \
V38=V38_part4+1.660555e+01*S40+2.166361e+01*S41 \
V39_part1=1.032811e+01*S0+1.000000e+04*S1+2.026242e+01*S2+1.000000e+04*S3+0.000000e+00*S4+2.044820e+01*S5+3.792265e+02*S6+(-1.108494e+02)*S7+(-1.977865e+00)*S8+7.180130e-01*S9 \
V39_part2=V39_part1+7.064182e+03*S10+6.515814e+00*S11+1.754970e-02*S12+7.010870e+00*S13+5.744304e+00*S14+6.349460e+00*S15+5.739539e+00*S16+3.966813e+00*S17+2.519697e+01*S18+6.613604e+00*S19 \
V39_part3=V39_part2+3.376491e+02*S20+1.064917e+01*S21+1.000000e+04*S22+5.437157e+02*S23+7.638135e+00*S24+5.974451e+01*S25+1.000000e+04*S26+1.000000e+04*S27+8.729158e+00*S28+2.386426e+00*S29 \
V39_part4=V39_part3+7.659774e+00*S30+3.375813e+01*S31+7.938970e+00*S32+6.365077e+01*S33+5.243279e+00*S34+6.448933e+00*S35+4.427886e+00*S36+3.385461e+00*S37+8.052841e+00*S38+(-3.527831e+02)*S39 \
V39=V39_part4+2.361640e+01*S40+2.504635e+00*S41 \
V40_part1=(-7.038472e+00)*S0+8.929972e+03*S1+(-2.015501e+01)*S2+(-5.208624e+03)*S3+0.000000e+00*S4+(-3.607374e+00)*S5+(-1.492025e+02)*S6+7.746047e+01*S7+2.263261e+00*S8+(-8.352298e-01)*S9 \
V40_part2=V40_part1+(-1.706652e+03)*S10+(-2.920883e+00)*S11+(-1.067715e+00)*S12+(-6.238097e-01)*S13+(-1.158203e+00)*S14+(-5.218181e+00)*S15+(-1.256571e+00)*S16+(-2.692971e+00)*S17+(-1.212685e+01)*S18+(-2.329841e+00)*S19 \
V40_part3=V40_part2+(-1.102427e+00)*S20+1.204822e+00*S21+1.000000e+04*S22+(-1.124598e+01)*S23+(-8.073286e+00)*S24+5.454939e+01*S25+1.000000e+04*S26+(-5.205599e+01)*S27+(-5.798854e+00)*S28+(-1.069930e+00)*S29 \
V40_part4=V40_part3+(-7.832030e+00)*S30+(-3.987342e+00)*S31+(-1.269835e+00)*S32+(-4.830273e+01)*S33+(-4.110381e+00)*S34+(-3.636390e+00)*S35+(-3.144556e+00)*S36+(-1.664417e+00)*S37+(-2.761723e+00)*S38+(-2.949473e+03)*S39 \
V40=V40_part4+(-3.808424e+00)*S40+(-9.666597e-01)*S41 \
V41_part1=(-4.313131e+00)*S0+(-1.000000e+04)*S1+1.351477e+00*S2+(-6.583476e+03)*S3+0.000000e+00*S4+(-1.413727e+01)*S5+(-1.577980e+02)*S6+2.714631e+02*S7+8.370301e+00*S8+2.568693e-01*S9 \
V41_part2=V41_part1+(-9.605124e+03)*S10+(-2.464086e+00)*S11+1.872931e+01*S12+(-6.203422e+00)*S13+(-3.878184e+00)*S14+4.927794e-02*S15+(-4.254317e+00)*S16+8.885272e-01*S17+(-2.646437e+01)*S18+(-2.951710e+00)*S19 \
V41_part3=V41_part2+(-6.178714e+02)*S20+(-1.527412e+01)*S21+9.108210e+03*S22+(-9.888799e+02)*S23+(-2.613931e+00)*S24+3.941391e+02*S25+1.000000e+04*S26+(-5.738863e-03)*S27+(-4.423781e+00)*S28+(-7.756519e-01)*S29 \
V41_part4=V41_part3+(-2.625265e+00)*S30+(-4.726938e+01)*S31+(-8.411207e+00)*S32+4.143911e+03*S33+1.042307e-01*S34+(-3.074568e-02)*S35+(-2.784362e+00)*S36+(-1.712172e+00)*S37+(-5.177480e+00)*S38+8.456839e+03*S39 \
V41=V41_part4+(-3.193067e+01)*S40+(-1.259623e+00)*S41 \
V42_part1=0.000000e+00*S0+3.975676e+00*S1+(-1.994151e+00)*S2+4.452210e+00*S3+0.000000e+00*S4+0.000000e+00*S5+2.021135e+01*S6+1.351551e+01*S7+7.250873e-02*S8+0.000000e+00*S9 \
V42_part2=V42_part1+0.000000e+00*S10+0.000000e+00*S11+3.519342e+01*S12+0.000000e+00*S13+0.000000e+00*S14+8.962287e+00*S15+0.000000e+00*S16+1.153029e+00*S17+0.000000e+00*S18+4.146129e+01*S19 \
V42_part3=V42_part2+0.000000e+00*S20+0.000000e+00*S21+(-2.839957e+00)*S22+(-8.334363e+00)*S23+1.201719e+01*S24+(-2.040765e+01)*S25+0.000000e+00*S26+1.425667e+01*S27+(-1.236487e+01)*S28+0.000000e+00*S29 \
V42_part4=V42_part3+3.743954e-01*S30+0.000000e+00*S31+0.000000e+00*S32+2.863473e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+(-2.460102e-01)*S37+(-6.054353e+01)*S38+0.000000e+00*S39 \
V42=V42_part4+0.000000e+00*S40+0.000000e+00*S41 \
V43_part1=0.000000e+00*S0+6.345238e+01*S1+6.573688e+01*S2+3.402457e+01*S3+0.000000e+00*S4+0.000000e+00*S5+8.405153e+01*S6+4.874259e-01*S7+6.249763e+01*S8+0.000000e+00*S9 \
V43_part2=V43_part1+0.000000e+00*S10+0.000000e+00*S11+6.181663e+01*S12+0.000000e+00*S13+0.000000e+00*S14+5.175779e+01*S15+0.000000e+00*S16+6.743712e+01*S17+0.000000e+00*S18+8.937751e+01*S19 \
V43_part3=V43_part2+0.000000e+00*S20+0.000000e+00*S21+5.663428e+01*S22+2.090521e+02*S23+5.169210e+01*S24+5.745024e+01*S25+0.000000e+00*S26+(-2.617091e+01)*S27+4.819107e+01*S28+0.000000e+00*S29 \
V43_part4=V43_part3+4.826362e+01*S30+0.000000e+00*S31+0.000000e+00*S32+4.129014e+01*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+(-1.287110e+01)*S37+7.482406e+01*S38+0.000000e+00*S39 \
V43=V43_part4+0.000000e+00*S40+0.000000e+00*S41 \
V44_part1=0.000000e+00*S0+1.112446e+01*S1+3.373023e+01*S2+1.467708e+01*S3+0.000000e+00*S4+0.000000e+00*S5+(-3.484628e+00)*S6+(-4.181949e-02)*S7+(-1.808743e+00)*S8+0.000000e+00*S9 \
V44_part2=V44_part1+0.000000e+00*S10+0.000000e+00*S11+1.606209e+01*S12+0.000000e+00*S13+0.000000e+00*S14+7.892004e+00*S15+0.000000e+00*S16+1.866993e+01*S17+0.000000e+00*S18+(-6.144445e+00)*S19 \
V44_part3=V44_part2+0.000000e+00*S20+0.000000e+00*S21+5.384646e+01*S22+(-1.885648e+02)*S23+3.291731e+01*S24+2.052390e+01*S25+0.000000e+00*S26+2.857434e+01*S27+6.034018e+01*S28+0.000000e+00*S29 \
V44_part4=V44_part3+5.023058e+01*S30+0.000000e+00*S31+0.000000e+00*S32+4.241898e+01*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+1.149393e+02*S37+5.944688e+01*S38+0.000000e+00*S39 \
V44=V44_part4+0.000000e+00*S40+0.000000e+00*S41 \
V45_part1=2.957583e+01*S0+1.838640e+03*S1+4.013571e+01*S2+(-1.999294e+03)*S3+5.189520e+00*S4+1.000000e+04*S5+2.069341e+01*S6+(-3.780457e+02)*S7+(-4.833351e+00)*S8+8.294555e+01*S9 \
V45_part2=V45_part1+1.413540e+03*S10+(-1.999258e+03)*S11+7.175111e-01*S12+3.490226e+00*S13+(-2.470992e+01)*S14+3.583104e+01*S15+(-3.450897e+01)*S16+4.486974e+01*S17+2.405120e+00*S18+(-4.389355e+00)*S19 \
V45_part3=V45_part2+(-3.717869e-03)*S20+3.378937e+00*S21+1.038976e+00*S22+(-6.550951e+02)*S23+4.199037e+01*S24+9.186617e-01*S25+3.563548e+00*S26+(-6.331059e+00)*S27+2.278575e+01*S28+2.069474e+01*S29 \
V45_part4=V45_part3+3.275538e+01*S30+1.053038e+00*S31+1.415040e+02*S32+2.677185e+01*S33+2.108969e+01*S34+1.039815e+01*S35+1.000000e+04*S36+1.273388e+03*S37+2.522309e+00*S38+3.554187e+01*S39 \
V45=V45_part4+(-3.609534e+00)*S40+1.643732e+01*S41 \
V46_part1=1.073286e-01*S0+7.032932e+02*S1+1.276095e+01*S2+(-5.267323e-01)*S3+(-1.147852e+00)*S4+1.181518e+02*S5+(-7.576068e+00)*S6+2.690420e+02*S7+(-1.188538e+01)*S8+(-4.431912e+01)*S9 \
V46_part2=V46_part1+(-4.626483e+03)*S10+(-7.617361e-01)*S11+1.003840e+00*S12+3.662132e+00*S13+3.377212e+02*S14+1.025344e+02*S15+(-4.897884e-01)*S16+1.047308e+01*S17+5.245658e-01*S18+(-1.647361e+00)*S19 \
V46_part3=V46_part2+(-1.945533e+00)*S20+3.954363e+00*S21+(-1.656502e+00)*S22+(-7.417568e-01)*S23+2.908184e+01*S24+(-2.650727e-01)*S25+2.332500e+00*S26+4.504937e+01*S27+4.521421e+01*S28+1.366419e-01*S29 \
V46_part4=V46_part3+1.974461e+01*S30+(-1.347064e+00)*S31+6.853637e+00*S32+1.587938e+01*S33+(-3.368400e+01)*S34+3.785854e+00*S35+1.000000e+04*S36+(-6.089162e+02)*S37+(-1.823149e+00)*S38+8.122928e+01*S39 \
V46=V46_part4+(-3.809779e-03)*S40+5.376112e+00*S41 \
V47_part1=(-3.127914e+01)*S0+1.000000e+04*S1+(-3.157840e+01)*S2+1.000000e+04*S3+(-2.265182e+00)*S4+1.000000e+04*S5+(-1.458604e+01)*S6+7.492939e+02*S7+8.677197e+01*S8+(-5.588089e+00)*S9 \
V47_part2=V47_part1+3.214686e+03*S10+1.000000e+04*S11+2.244748e-01*S12+(-4.296998e+00)*S13+(-1.368694e+02)*S14+(-5.790681e+01)*S15+1.759572e+02*S16+(-3.814606e+01)*S17+(-1.668960e+00)*S18+2.961937e+01*S19 \
V47_part3=V47_part2+1.344750e+01*S20+(-6.437736e+00)*S21+3.171842e+00*S22+3.281107e+03*S23+(-8.820972e+01)*S24+(-1.555904e-01)*S25+(-9.007115e+00)*S26+(-1.482607e+00)*S27+(-7.631028e+01)*S28+(-3.538965e+01)*S29 \
V47_part4=V47_part3+(-6.737959e+01)*S30+1.667854e+00*S31+(-2.717948e+02)*S32+(-5.396921e+01)*S33+2.996392e+01*S34+(-2.342912e+01)*S35+1.000000e+04*S36+(-1.498801e+03)*S37+1.878794e+00*S38+(-1.057885e+02)*S39 \
V47=V47_part4+2.375058e+01*S40+(-3.523628e+01)*S41 \
V48_part1=(-3.566372e-01)*S0+0.000000e+00*S1+(-3.792115e-01)*S2+(-3.001705e-01)*S3+(-2.275049e-01)*S4+0.000000e+00*S5+(-1.408316e-01)*S6+(-1.304064e-01)*S7+0.000000e+00*S8+2.596202e-02*S9 \
V48_part2=V48_part1+(-3.799801e-01)*S10+0.000000e+00*S11+5.248625e-01*S12+(-1.369291e-01)*S13+0.000000e+00*S14+0.000000e+00*S15+(-8.114884e-01)*S16+0.000000e+00*S17+2.757070e-01*S18+(-4.609412e-01)*S19 \
V48_part3=V48_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+(-3.322964e-01)*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+(-3.328376e-02)*S27+0.000000e+00*S28+(-6.895291e-01)*S29 \
V48_part4=V48_part3+(-5.970622e-02)*S30+(-8.819791e-01)*S31+(-3.505653e-01)*S32+0.000000e+00*S33+(-4.216330e-01)*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+(-2.717782e+00)*S38+0.000000e+00*S39 \
V48=V48_part4+(-5.510386e-01)*S40+(-9.066139e-01)*S41 \
V49_part1=1.339699e+00*S0+0.000000e+00*S1+8.567048e-01*S2+7.287052e-01*S3+6.657083e-01*S4+0.000000e+00*S5+2.558613e-01*S6+4.344103e-01*S7+0.000000e+00*S8+1.638793e-01*S9 \
V49_part2=V49_part1+1.853198e+00*S10+0.000000e+00*S11+(-2.799405e-01)*S12+1.470174e+00*S13+0.000000e+00*S14+0.000000e+00*S15+1.361158e+00*S16+0.000000e+00*S17+2.123988e+00*S18+2.405507e+00*S19 \
V49_part3=V49_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+1.505790e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+1.571346e+00*S27+0.000000e+00*S28+3.990725e+00*S29 \
V49_part4=V49_part3+7.095459e-01*S30+7.907650e-01*S31+4.115839e+00*S32+0.000000e+00*S33+1.083982e+00*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+2.945893e+00*S38+0.000000e+00*S39 \
V49=V49_part4+2.129253e+00*S40+3.532509e+00*S41 \
V50_part1=4.226898e-01*S0+0.000000e+00*S1+3.310621e-01*S2+2.813102e-01*S3+9.250978e-01*S4+0.000000e+00*S5+5.001021e-01*S6+1.619874e-01*S7+0.000000e+00*S8+1.906142e-01*S9 \
V50_part2=V50_part1+6.380278e-01*S10+0.000000e+00*S11+(-3.261495e-01)*S12+3.794260e-01*S13+0.000000e+00*S14+0.000000e+00*S15+1.335515e+00*S16+0.000000e+00*S17+(-1.342617e-01)*S18+1.158467e+00*S19 \
V50_part3=V50_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+4.162014e-01*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+1.164424e-01*S27+0.000000e+00*S28+(-3.347328e+00)*S29 \
V50_part4=V50_part3+1.486464e-01*S30+6.202505e+00*S31+(-2.712191e+00)*S32+0.000000e+00*S33+8.346685e-02*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+2.982438e+00*S38+0.000000e+00*S39 \
V50=V50_part4+1.839987e+00*S40+(-8.388909e-01)*S41 \
V51_part1=1.420024e+01*S0+1.000000e+04*S1+2.783026e-01*S2+(-1.488369e+02)*S3+9.595593e+00*S4+(-2.643628e+02)*S5+0.000000e+00*S6+(-3.423705e+01)*S7+2.336845e+00*S8+7.916396e+00*S9 \
V51_part2=V51_part1+7.964241e+00*S10+8.310703e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+(-3.300666e+03)*S15+0.000000e+00*S16+(-5.632974e+02)*S17+(-1.248503e+02)*S18+0.000000e+00*S19 \
V51_part3=V51_part2+9.710519e+03*S20+5.546266e+02*S21+1.124133e+03*S22+(-9.605101e-01)*S23+8.209916e+00*S24+1.019026e+02*S25+5.848805e-01*S26+1.313212e+00*S27+(-2.565449e+00)*S28+0.000000e+00*S29 \
V51_part4=V51_part3+1.806184e+01*S30+4.865681e+01*S31+0.000000e+00*S32+(-2.330338e-01)*S33+1.285692e+02*S34+(-1.661099e+02)*S35+(-3.556174e+01)*S36+3.204096e+02*S37+2.240246e+02*S38+(-2.004946e+03)*S39 \
V51=V51_part4+0.000000e+00*S40+1.965297e+02*S41 \
V52_part1=3.394337e-01*S0+8.078340e+03*S1+(-8.684496e-01)*S2+3.295354e+02*S3+(-1.037204e+00)*S4+1.872170e+03*S5+0.000000e+00*S6+1.460712e+02*S7+3.398572e-01*S8+1.912939e+00*S9 \
V52_part2=V52_part1+(-1.908821e+00)*S10+1.611671e+01*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+(-8.458107e+01)*S15+0.000000e+00*S16+(-3.099060e+01)*S17+(-2.191185e+00)*S18+0.000000e+00*S19 \
V52_part3=V52_part2+9.710519e+03*S20+(-1.780021e+03)*S21+1.155142e+03*S22+(-7.220450e-01)*S23+(-2.025999e+02)*S24+(-1.508537e+01)*S25+(-5.010432e-01)*S26+(-4.228332e+00)*S27+(-3.383525e+00)*S28+0.000000e+00*S29 \
V52_part4=V52_part3+(-5.999115e+01)*S30+9.174746e+00*S31+0.000000e+00*S32+(-2.622060e+01)*S33+3.691098e+00*S34+2.419512e+02*S35+(-2.691025e+00)*S36+1.345457e+02*S37+(-2.242900e+02)*S38+3.228388e+02*S39 \
V52=V52_part4+0.000000e+00*S40+5.153928e+02*S41 \
V53_part1=(-1.322785e+01)*S0+(-1.000000e+04)*S1+8.968785e-01*S2+(-5.388398e+01)*S3+(-5.476655e+00)*S4+(-4.271950e+02)*S5+0.000000e+00*S6+(-8.367758e+00)*S7+(-2.949057e+00)*S8+(-5.681992e+00)*S9 \
V53_part2=V53_part1+(-9.044495e+00)*S10+(-2.911232e+01)*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+8.437621e+03*S15+0.000000e+00*S16+1.487216e+03*S17+6.311649e+02*S18+0.000000e+00*S19 \
V53_part3=V53_part2+(-3.853020e+01)*S20+1.370949e+03*S21+(-3.035510e+03)*S22+1.071103e+01*S23+4.292665e+02*S24+(-1.496058e+02)*S25+8.126110e-01*S26+6.507231e+00*S27+2.941996e+01*S28+0.000000e+00*S29 \
V53_part4=V53_part3+5.804274e+01*S30+1.116478e+02*S31+0.000000e+00*S32+7.324141e+01*S33+(-2.396612e+02)*S34+2.201308e+02*S35+1.885694e+03*S36+5.735364e+02*S37+3.468065e+02*S38+9.899862e+03*S39 \
V53=V53_part4+0.000000e+00*S40+1.071127e+03*S41 \
V54_part1=0.000000e+00*S0+0.000000e+00*S1+6.764185e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+(-1.256710e+00)*S8+0.000000e+00*S9 \
V54_part2=V54_part1+0.000000e+00*S10+6.466468e+00*S11+3.198097e+01*S12+0.000000e+00*S13+0.000000e+00*S14+(-1.489283e-01)*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V54_part3=V54_part2+(-3.563902e+02)*S20+3.013558e-01*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+6.615903e-01*S27+3.498150e-02*S28+0.000000e+00*S29 \
V54_part4=V54_part3+0.000000e+00*S30+0.000000e+00*S31+(-5.854221e-01)*S32+(-3.141472e-02)*S33+0.000000e+00*S34+0.000000e+00*S35+1.270586e-02*S36+(-4.810748e-01)*S37+0.000000e+00*S38+0.000000e+00*S39 \
V54=V54_part4+0.000000e+00*S40+(-3.140910e+03)*S41 \
V55_part1=0.000000e+00*S0+0.000000e+00*S1+(-8.362421e+00)*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+1.937471e+00*S8+0.000000e+00*S9 \
V55_part2=V55_part1+0.000000e+00*S10+(-4.237904e+00)*S11+6.082531e+00*S12+0.000000e+00*S13+0.000000e+00*S14+2.170435e-01*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V55_part3=V55_part2+(-8.039298e+02)*S20+4.809068e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+(-5.360477e-01)*S27+7.701028e-01*S28+0.000000e+00*S29 \
V55_part4=V55_part3+0.000000e+00*S30+0.000000e+00*S31+2.468469e+01*S32+6.646937e-01*S33+0.000000e+00*S34+0.000000e+00*S35+2.278270e+00*S36+2.209654e+00*S37+0.000000e+00*S38+0.000000e+00*S39 \
V55=V55_part4+0.000000e+00*S40+9.837207e+03*S41 \
V56_part1=0.000000e+00*S0+0.000000e+00*S1+7.629907e-01*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+1.555455e+00*S8+0.000000e+00*S9 \
V56_part2=V56_part1+0.000000e+00*S10+(-3.658298e+00)*S11+(-3.237115e+01)*S12+0.000000e+00*S13+0.000000e+00*S14+1.766109e-01*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V56_part3=V56_part2+5.894455e+03*S20+1.228228e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+(-5.262837e-01)*S27+(-2.070745e-01)*S28+0.000000e+00*S29 \
V56_part4=V56_part3+0.000000e+00*S30+0.000000e+00*S31+2.520933e+02*S32+1.899131e-02*S33+0.000000e+00*S34+0.000000e+00*S35+4.345574e+00*S36+1.553789e+00*S37+0.000000e+00*S38+0.000000e+00*S39 \
V56=V56_part4+0.000000e+00*S40+7.922716e+03*S41 \
V57_part1=0.000000e+00*S0+4.001488e-01*S1+6.208800e+03*S2+(-9.735421e-02)*S3+7.440045e+00*S4+0.000000e+00*S5+4.839591e+00*S6+0.000000e+00*S7+(-3.531289e-01)*S8+(-5.502093e+00)*S9 \
V57_part2=V57_part1+0.000000e+00*S10+2.292499e+00*S11+1.275057e+01*S12+(-2.077000e+01)*S13+(-1.999290e+03)*S14+0.000000e+00*S15+6.440014e+00*S16+8.829975e+00*S17+0.000000e+00*S18+6.037948e+00*S19 \
V57_part3=V57_part2+1.383374e+02*S20+5.950123e+00*S21+0.000000e+00*S22+2.015164e+00*S23+8.604213e+00*S24+9.002145e+00*S25+0.000000e+00*S26+1.787380e+03*S27+0.000000e+00*S28+9.945173e-01*S29 \
V57_part4=V57_part3+0.000000e+00*S30+2.426807e-01*S31+1.144009e+00*S32+0.000000e+00*S33+0.000000e+00*S34+1.614984e+02*S35+0.000000e+00*S36+8.021145e+01*S37+3.503448e+02*S38+2.911656e+00*S39 \
V57=V57_part4+3.430267e+01*S40+1.513825e+00*S41 \
V58_part1=0.000000e+00*S0+(-1.006805e-01)*S1+(-8.303294e+03)*S2+1.739774e+00*S3+2.098943e+00*S4+0.000000e+00*S5+4.131831e+00*S6+0.000000e+00*S7+6.108292e-01*S8+1.169953e+01*S9 \
V58_part2=V58_part1+0.000000e+00*S10+(-1.289851e+00)*S11+2.367844e+00*S12+(-1.431933e+00)*S13+(-6.865047e-01)*S14+0.000000e+00*S15+3.733437e+00*S16+1.475062e+02*S17+0.000000e+00*S18+4.655627e+00*S19 \
V58_part3=V58_part2+3.853316e+00*S20+(-1.355344e+01)*S21+0.000000e+00*S22+7.630229e+00*S23+(-1.946996e+01)*S24+(-7.773255e+00)*S25+0.000000e+00*S26+3.352825e+00*S27+0.000000e+00*S28+(-1.462695e+00)*S29 \
V58_part4=V58_part3+0.000000e+00*S30+(-4.313719e-01)*S31+(-1.293587e+00)*S32+0.000000e+00*S33+0.000000e+00*S34+1.903993e+01*S35+0.000000e+00*S36+6.068219e+01*S37+1.729456e+00*S38+(-2.404144e+00)*S39 \
V58=V58_part4+2.235382e+01*S40+(-1.938043e+00)*S41 \
V59_part1=0.000000e+00*S0+(-1.084645e-01)*S1+2.353896e+03*S2+(-1.369682e+00)*S3+(-4.220136e+00)*S4+0.000000e+00*S5+(-7.006704e+00)*S6+0.000000e+00*S7+(-1.089379e-01)*S8+5.566818e+00*S9 \
V59_part2=V59_part1+0.000000e+00*S10+(-1.916379e+00)*S11+(-2.491436e+01)*S12+1.078397e+02*S13+1.000000e+04*S14+0.000000e+00*S15+(-1.023575e+01)*S16+1.155906e+01*S17+0.000000e+00*S18+(-1.361909e+01)*S19 \
V59_part3=V59_part2+(-2.615852e+02)*S20+1.181709e+00*S21+0.000000e+00*S22+(-1.267897e+01)*S23+8.149332e+00*S24+(-7.742839e-01)*S25+0.000000e+00*S26+2.593803e+00*S27+0.000000e+00*S28+4.496729e+00*S29 \
V59_part4=V59_part3+0.000000e+00*S30+7.744143e+00*S31+2.284841e+00*S32+0.000000e+00*S33+0.000000e+00*S34+2.891670e+03*S35+0.000000e+00*S36+2.120763e+03*S37+1.901673e+01*S38+(-8.217598e-02)*S39 \
V59=V59_part4+(-5.688807e+01)*S40+4.950844e+00*S41 \
V60_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+6.412445e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V60_part2=V60_part1+0.000000e+00*S10+(-7.658182e-01)*S11+(-3.116305e-02)*S12+0.000000e+00*S13+(-2.855307e-01)*S14+5.736403e+01*S15+0.000000e+00*S16+3.532043e+00*S17+1.242188e+03*S18+0.000000e+00*S19 \
V60_part3=V60_part2+(-5.376781e-01)*S20+(-9.627405e-01)*S21+0.000000e+00*S22+0.000000e+00*S23+(-1.575252e+01)*S24+0.000000e+00*S25+0.000000e+00*S26+4.232718e-01*S27+0.000000e+00*S28+0.000000e+00*S29 \
V60_part4=V60_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+(-9.312063e-01)*S33+0.000000e+00*S34+(-1.447873e-02)*S35+0.000000e+00*S36+(-1.853545e+01)*S37+0.000000e+00*S38+0.000000e+00*S39 \
V60=V60_part4+0.000000e+00*S40+0.000000e+00*S41 \
V61_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+9.095159e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V61_part2=V61_part1+0.000000e+00*S10+2.248277e+00*S11+1.729896e+00*S12+0.000000e+00*S13+6.564487e-01*S14+5.849738e+01*S15+0.000000e+00*S16+1.646506e+00*S17+1.000000e+04*S18+0.000000e+00*S19 \
V61_part3=V61_part2+2.036723e+00*S20+6.518272e+00*S21+0.000000e+00*S22+0.000000e+00*S23+1.746698e+01*S24+0.000000e+00*S25+0.000000e+00*S26+1.025664e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V61_part4=V61_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+2.736571e+01*S33+0.000000e+00*S34+6.571587e-01*S35+0.000000e+00*S36+3.904119e+03*S37+0.000000e+00*S38+0.000000e+00*S39 \
V61=V61_part4+0.000000e+00*S40+0.000000e+00*S41 \
V62_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+8.842000e+01*S7+0.000000e+00*S8+0.000000e+00*S9 \
V62_part2=V62_part1+0.000000e+00*S10+2.054814e+00*S11+(-6.472534e-01)*S12+0.000000e+00*S13+3.734876e-01*S14+1.721057e+02*S15+0.000000e+00*S16+2.106343e+02*S17+1.000000e+04*S18+0.000000e+00*S19 \
V62_part3=V62_part2+(-4.677948e-01)*S20+8.396335e-01*S21+0.000000e+00*S22+0.000000e+00*S23+6.476430e+01*S24+0.000000e+00*S25+0.000000e+00*S26+4.480992e-02*S27+0.000000e+00*S28+0.000000e+00*S29 \
V62_part4=V62_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+(-1.060457e+00)*S33+0.000000e+00*S34+(-5.911740e-01)*S35+0.000000e+00*S36+4.495738e+03*S37+0.000000e+00*S38+0.000000e+00*S39 \
V62=V62_part4+0.000000e+00*S40+0.000000e+00*S41 \
_P0=V0+V1*radius_+V2*w_ \
_P1=0.5*(_P0+sqrt(_P0*_P0+0.001)) \
_P2=1e-15*_P1 \
_P3=V3+V4*radius_+V5/w_ \
_P4=0.5*(_P3+sqrt(_P3*_P3+0.001)) \
_P5=V6+V7*radius_+V8*w_ \
_P6=0.5*(_P5+sqrt(_P5*_P5+0.001)) \
_P7=1e-09*_P6 \
_P8=1e-09*_P6 \
_P9=V9+V10*radius_+V11/w_ \
_P10=0.5*(_P9+sqrt(_P9*_P9+0.001)) \
_P11=V12+V13*radius_+V14*w_ \
_P12=0.5*(_P11+sqrt(_P11*_P11+0.001)) \
_P13=1e-09*_P12 \
_P14=V15+V16*radius_+V17*w_ \
_P15=0.5*(atan(2*_P14)/1.5708+1) \
_P16=0.7064*_P15 \
_P17=0.7064*_P15 \
_P18=V18+V19*radius_+V20*w_ \
_P19=0.5*(_P18+sqrt(_P18*_P18+0.001)) \
_P20=V21+V22*radius_+V23*w_ \
_P21=0.5*(_P20+sqrt(_P20*_P20+0.001)) \
_P22=V24+V25*radius_+V26*w_ \
_P23=0.5*(_P22+sqrt(_P22*_P22+0.001)) \
_P24=V27+V28*radius_+V29*w_ \
_P25=0.5*(_P24+sqrt(_P24*_P24+0.001)) \
_P26=V30+V31*radius_+V32*w_ \
_P27=0.5*(_P26+sqrt(_P26*_P26+0.001)) \
_P28=V33+V34*radius_+V35*w_ \
_P29=0.5*(_P28+sqrt(_P28*_P28+0.001)) \
_P30=V36+V37*radius_+V38*w_ \
_P31=0.5*(_P30+sqrt(_P30*_P30+0.001)) \
_P32=V39+V40*radius_+V41*w_ \
_P33=0.5*(_P32+sqrt(_P32*_P32+0.001)) \
_P34=V42+V43*radius_+V44*w_ \
_P35=0.5*(_P34+sqrt(_P34*_P34+0.001)) \
_P36=1e-14*_P19 \
_P37=100*_P21 \
_P38=1e-15*_P23 \
_P39=1e-14*_P25 \
_P40=100*_P27 \
_P41=1e-15*_P29 \
_P42=1e-14*_P31 \
_P43=100*_P33 \
_P44=1e-15*_P35 \
_P45=V45+V46*radius_+V47*w_ \
_P46=0.5*(_P45+sqrt(_P45*_P45+0.001)) \
_P47=V48+V49*radius_+V50*w_ \
_P48=0.5*(_P47+sqrt(_P47*_P47+0.001)) \
_P49=100*_P46 \
_P50=1e-13*_P48 \
_P51=V51+V52*radius_+V53*w_ \
_P52=0.5*(_P51+sqrt(_P51*_P51+0.001)) \
_P53=V54+V55*radius_+V56*w_ \
_P54=0.5*(_P53+sqrt(_P53*_P53+0.001)) \
_P55=100*_P52 \
_P56=1e-13*_P54 \
_P57=V57+V58*radius_+V59*w_ \
_P58=0.5*(_P57+sqrt(_P57*_P57+0.001)) \
_P59=V60+V61*radius_+V62*w_ \
_P60=0.5*(_P59+sqrt(_P59*_P59+0.001)) \
_P61=100*_P58 \
_P62=1e-13*_P60
cs (PLUS MINUS) capacitor c=_P2
rs1_1 (PLUS n1_1) resistor r=_P4*(1+drs_ind_rf_psub) tc1=0.003
ls1_1 (n1_1 ni_1) inductor l=_P7*(1+dls_ind_rf_psub)
rs2_1 (ni_1 n2_1) resistor r=_P4*(1+drs_ind_rf_psub) tc1=0.003
ls2_1 (n2_1 MINUS) inductor l=_P8*(1+dls_ind_rf_psub)
rs1_2 (PLUS n1_2) resistor r=_P10*(1+drs_ind_rf_psub) tc1=0.003
ls1_2 (n1_2 MINUS) inductor l=_P13*(1+dls_ind_rf_psub)
k1 mutual_inductor coupling=_P16 ind1=ls1_1 ind2=ls1_2
k2 mutual_inductor coupling=_P17 ind1=ls2_1 ind2=ls1_2
c_1_sub (PLUS _n1_1_sub) capacitor c=_P36
rs_1_sub (_n1_1_sub PSUB) resistor r=_P37
cs_1_sub (_n1_1_sub PSUB) capacitor c=_P38
c_2_sub (MINUS _n1_2_sub) capacitor c=_P39
rs_2_sub (_n1_2_sub PSUB) resistor r=_P40
cs_2_sub (_n1_2_sub PSUB) capacitor c=_P41
c_3_sub (ni_1 _n1_3_sub) capacitor c=_P42
rs_3_sub (_n1_3_sub PSUB) resistor r=_P43
cs_3_sub (_n1_3_sub PSUB) capacitor c=_P44
rx_1_2_sub (_n1_1_sub _n1_2_sub) resistor r=_P49
cx_1_2_sub (_n1_1_sub _n1_2_sub) capacitor c=_P50
rx_1_3_sub (_n1_1_sub _n1_3_sub) resistor r=_P55
cx_1_3_sub (_n1_1_sub _n1_3_sub) capacitor c=_P56
rx_2_3_sub (_n1_2_sub _n1_3_sub) resistor r=_P61
cx_2_3_sub (_n1_2_sub _n1_3_sub) capacitor c=_P62
ends ind_rf_psub
