`timescale 1ns / 1ns

module simu_top();

   reg clk;//system input
   reg wen;//system input
   reg wbuf;//system input
   reg cal;//system input
   reg [8:0] addra;//system input
   reg [15:0]dina;//sys input and CIM input
   wire cal_done;//system output
   wire [7:0] douta; //system output

   reg clk_CIM_a;
   wire clk_CIM;// CIM input
   wire [15:0]q_in_cim;//CIM output
   wire comp;//CIM input
   wire model;//CIM input
   wire wait_;//CIM input
   wire inbit;//CIM input
   wire set;//CIM input
   wire read;//CIM input
   wire [8:0]a;//CIM input
   wire wrt;//CIM input
   wire wrtbuf;//CIM input

   
   wire [3:0]cim_a;
   wire cal_b; 

    
    real    CLK_PEROID = 100;
    real    HIGH_RATE = 0.4;
    always begin
        clk = 1 ; #(CLK_PEROID*0.5) ;
        clk = 0 ; #(CLK_PEROID*0.5) ;
    end
    always begin
        clk_CIM_a = 1 ; #(CLK_PEROID*HIGH_RATE) ;
        clk_CIM_a = 0 ; #(CLK_PEROID*(1-HIGH_RATE));
    end

    assign #(CLK_PEROID*(0.5-HIGH_RATE)*0.5) clk_CIM = clk_CIM_a;

    IOw iow(
     .clk(clk),
     .wen(wen),
     .wbuf(wbuf),
     .cal(cal),
     .a_in(addra),
     .cim_a(cim_a),
     .read(read),
     .a_out(a),
     .wrt(wrt), 
     .wrtbuf(wrtbuf),
     .cal_b(cal_b)//cal_b�źŲ���״̬���Ŀ���
    );

   wire [7:0]SMw_data;
   SMw smw(
    .clk(clk),
    .cal_b(cal_b),
    .q(q_in_cim),
    .cim_a(cim_a),
    .a(addra[4:0]),//adderess of out ,form system IO
    .comp(comp),
    .model(model),
    .wait_(wait_),
    .inbit(inbit),
    .set(set),
    .read(read),
    .cal_done(cal_done),
    .data_out(SMw_data)
    );
    reg eact;//system input
    ACT act(
        .eact(eact),
        .data_in(SMw_data),
        .data_out(douta)
        );
        
    SRAM_CIM dut(
        .a(a), 
        .d(dina),
        .q(q_in_cim),
        .clk(clk_CIM),
        .comp(comp),
        .inbit(inbit),
        .model(model),
        .read(read),
        .set(set),
        .wait_(wait_),
        .wrt(wrt),
        .wrtbuf(wrtbuf)
    );
   //task define
    task test_writeBUF;
        input [4:0] B_addr;
        input [15:0] B_data;

        begin
            addra[4:0] = B_addr;
            dina = ~B_data;
            wen = 1'b1;
            wbuf = 1'b1;
            #(CLK_PEROID)
            wen = 1'b0;
            wbuf = 1'b0;
            #(CLK_PEROID);
        end
    endtask


    task test_writeARY;
        input [8:0] A_addr;
        input [15:0] A_data;

        begin
            addra = A_addr;
            dina = ~A_data;
            wen = 1'b1;
            wbuf = 1'b0;
            #(CLK_PEROID)
            wen = 1'b0; 
            wbuf = 1'b0;
            #(CLK_PEROID);
        end
    endtask

    task test_cal;
        begin
            cal = 1'b1;
            #(CLK_PEROID *30) cal = 1'b0;
            #(CLK_PEROID);
        end
    endtask

    task test_read;
        input[4:0] R_addr;
        input is_ACT;
        reg [7:0]R_data;
        begin   
            addra[4:0] = R_addr;
            eact = is_ACT;
            R_data = douta;
            $display("cALCULATION Result is %d",R_data);
        end
    endtask
   //
    initial begin
        # (CLK_PEROID /  2);
        addra = 9'b0;//system input
        dina = 16'b0;//sys input
        wen = 1'b0;//sys input
        wbuf = 1'b0;//sys input
        cal = 1'b0;//sys input
        eact = 1'b0;//sys input
		$fsdbDumpfile("vcs_simutop.fsdb");
		$fsdbDumpvars;
        $fsdbDumpMDA();
    //writeBUF
        test_writeBUF(5'd0,16'b1111111111111111);
        test_writeBUF(5'd1,16'b1111111111111111);
        test_writeBUF(5'd2,16'b1111111111111111);
        test_writeBUF(5'd3,16'b1111111111111111);
        test_writeBUF(5'd4,16'b1111111111111111);
        test_writeBUF(5'd5,16'b1111111111111111);
        test_writeBUF(5'd6,16'b1111111111111111);
        test_writeBUF(5'd7,16'b1111111111111111);
        test_writeBUF(5'd8,16'b1111111111111111);
        test_writeBUF(5'd9,16'b1111111111111111);
        test_writeBUF(5'd10,16'b1111111111111111);
        test_writeBUF(5'd11,16'b1111111111111111);
        test_writeBUF(5'd12,16'b1111111111111111);
        test_writeBUF(5'd13,16'b1111111111111111);
        test_writeBUF(5'd14,16'b1111111111111111);
        test_writeBUF(5'd15,16'b1111111111111111);
        test_writeBUF(5'd16,16'b1111111111111111);
        test_writeBUF(5'd17,16'b1111111111111111);
        test_writeBUF(5'd18,16'b1111111111111111);
        test_writeBUF(5'd19,16'b1111111111111111);
        test_writeBUF(5'd20,16'b1111111111111111);
        test_writeBUF(5'd21,16'b1111111111111111);
        test_writeBUF(5'd22,16'b1111111111111111);
        test_writeBUF(5'd23,16'b1111111111111111);
        test_writeBUF(5'd24,16'b1111111111111111);
        test_writeBUF(5'd25,16'b1111111111111111);
        test_writeBUF(5'd26,16'b1111111111111111);
        test_writeBUF(5'd27,16'b1111111111111111);
        test_writeBUF(5'd28,16'b1111111111111111);
        test_writeBUF(5'd29,16'b1111111111111111);
        test_writeBUF(5'd30,16'b1111111111111111);
        test_writeBUF(5'd31,16'b1111111111111111);
    //
    //writeARY
        test_writeARY(9'd0,16'b1010101010101010);
        test_writeARY(9'd1,16'b1010101010101010);
        test_writeARY(9'd2,16'b1010101010101010);
        test_writeARY(9'd3,16'b1010101010101010);
        test_writeARY(9'd4,16'b1010101010101010);
        test_writeARY(9'd5,16'b1010101010101010);
        test_writeARY(9'd6,16'b1010101010101010);
        test_writeARY(9'd7,16'b1010101010101010);
        test_writeARY(9'd8,16'b1010101010101010);
        test_writeARY(9'd9,16'b1010101010101010);
        test_writeARY(9'd10,16'b1010101010101010);
        test_writeARY(9'd11,16'b1010101010101010);
        test_writeARY(9'd12,16'b1010101010101010);
        test_writeARY(9'd13,16'b1010101010101010);
        test_writeARY(9'd14,16'b1010101010101010);
        test_writeARY(9'd15,16'b1010101010101010);
        test_writeARY(9'd16,16'b1010101010101010);
        test_writeARY(9'd17,16'b1010101010101010);
        test_writeARY(9'd18,16'b1010101010101010);
        test_writeARY(9'd19,16'b1010101010101010);
        test_writeARY(9'd20,16'b1010101010101010);
        test_writeARY(9'd21,16'b1010101010101010);
        test_writeARY(9'd22,16'b1010101010101010);
        test_writeARY(9'd23,16'b1010101010101010);
        test_writeARY(9'd24,16'b1010101010101010);
        test_writeARY(9'd25,16'b1010101010101010);
        test_writeARY(9'd26,16'b1010101010101010);
        test_writeARY(9'd27,16'b1010101010101010);
        test_writeARY(9'd28,16'b1010101010101010);
        test_writeARY(9'd29,16'b1010101010101010);
        test_writeARY(9'd30,16'b1010101010101010);
        test_writeARY(9'd31,16'b1010101010101010);
        test_writeARY(9'd32,16'b1010101010101010);
        test_writeARY(9'd33,16'b1010101010101010);
        test_writeARY(9'd34,16'b1010101010101010);
        test_writeARY(9'd35,16'b1010101010101010);
        test_writeARY(9'd36,16'b1010101010101010);
        test_writeARY(9'd37,16'b1010101010101010);
        test_writeARY(9'd38,16'b1010101010101010);
        test_writeARY(9'd39,16'b1010101010101010);
        test_writeARY(9'd40,16'b1010101010101010);
        test_writeARY(9'd41,16'b1010101010101010);
        test_writeARY(9'd42,16'b1010101010101010);
        test_writeARY(9'd43,16'b1010101010101010);
        test_writeARY(9'd44,16'b1010101010101010);
        test_writeARY(9'd45,16'b1010101010101010);
        test_writeARY(9'd46,16'b1010101010101010);
        test_writeARY(9'd47,16'b1010101010101010);
        test_writeARY(9'd48,16'b1010101010101010);
        test_writeARY(9'd49,16'b1010101010101010);
        test_writeARY(9'd50,16'b1010101010101010);
        test_writeARY(9'd51,16'b1010101010101010);
        test_writeARY(9'd52,16'b1010101010101010);
        test_writeARY(9'd53,16'b1010101010101010);
        test_writeARY(9'd54,16'b1010101010101010);
        test_writeARY(9'd55,16'b1010101010101010);
        test_writeARY(9'd56,16'b1010101010101010);
        test_writeARY(9'd57,16'b1010101010101010);
        test_writeARY(9'd58,16'b1010101010101010);
        test_writeARY(9'd59,16'b1010101010101010);
        test_writeARY(9'd60,16'b1010101010101010);
        test_writeARY(9'd61,16'b1010101010101010);
        test_writeARY(9'd62,16'b1010101010101010);
        test_writeARY(9'd63,16'b1010101010101010);
        test_writeARY(9'd64,16'b1010101010101010);
        test_writeARY(9'd65,16'b1010101010101010);
        test_writeARY(9'd66,16'b1010101010101010);
        test_writeARY(9'd67,16'b1010101010101010);
        test_writeARY(9'd68,16'b1010101010101010);
        test_writeARY(9'd69,16'b1010101010101010);
        test_writeARY(9'd70,16'b1010101010101010);
        test_writeARY(9'd71,16'b1010101010101010);
        test_writeARY(9'd72,16'b1010101010101010);
        test_writeARY(9'd73,16'b1010101010101010);
        test_writeARY(9'd74,16'b1010101010101010);
        test_writeARY(9'd75,16'b1010101010101010);
        test_writeARY(9'd76,16'b1010101010101010);
        test_writeARY(9'd77,16'b1010101010101010);
        test_writeARY(9'd78,16'b1010101010101010);
        test_writeARY(9'd79,16'b1010101010101010);
        test_writeARY(9'd80,16'b1010101010101010);
        test_writeARY(9'd81,16'b1010101010101010);
        test_writeARY(9'd82,16'b1010101010101010);
        test_writeARY(9'd83,16'b1010101010101010);
        test_writeARY(9'd84,16'b1010101010101010);
        test_writeARY(9'd85,16'b1010101010101010);
        test_writeARY(9'd86,16'b1010101010101010);
        test_writeARY(9'd87,16'b1010101010101010);
        test_writeARY(9'd88,16'b1010101010101010);
        test_writeARY(9'd89,16'b1010101010101010);
        test_writeARY(9'd90,16'b1010101010101010);
        test_writeARY(9'd91,16'b1010101010101010);
        test_writeARY(9'd92,16'b1010101010101010);
        test_writeARY(9'd93,16'b1010101010101010);
        test_writeARY(9'd94,16'b1010101010101010);
        test_writeARY(9'd95,16'b1010101010101010);
        test_writeARY(9'd96,16'b1010101010101010);
        test_writeARY(9'd97,16'b1010101010101010);
        test_writeARY(9'd98,16'b1010101010101010);
        test_writeARY(9'd99,16'b1010101010101010);
        test_writeARY(9'd100,16'b1010101010101010);
        test_writeARY(9'd101,16'b1010101010101010);
        test_writeARY(9'd102,16'b1010101010101010);
        test_writeARY(9'd103,16'b1010101010101010);
        test_writeARY(9'd104,16'b1010101010101010);
        test_writeARY(9'd105,16'b1010101010101010);
        test_writeARY(9'd106,16'b1010101010101010);
        test_writeARY(9'd107,16'b1010101010101010);
        test_writeARY(9'd108,16'b1010101010101010);
        test_writeARY(9'd109,16'b1010101010101010);
        test_writeARY(9'd110,16'b1010101010101010);
        test_writeARY(9'd111,16'b1010101010101010);
        test_writeARY(9'd112,16'b1010101010101010);
        test_writeARY(9'd113,16'b1010101010101010);
        test_writeARY(9'd114,16'b1010101010101010);
        test_writeARY(9'd115,16'b1010101010101010);
        test_writeARY(9'd116,16'b1010101010101010);
        test_writeARY(9'd117,16'b1010101010101010);
        test_writeARY(9'd118,16'b1010101010101010);
        test_writeARY(9'd119,16'b1010101010101010);
        test_writeARY(9'd120,16'b1010101010101010);
        test_writeARY(9'd121,16'b1010101010101010);
        test_writeARY(9'd122,16'b1010101010101010);
        test_writeARY(9'd123,16'b1010101010101010);
        test_writeARY(9'd124,16'b1010101010101010);
        test_writeARY(9'd125,16'b1010101010101010);
        test_writeARY(9'd126,16'b1010101010101010);
        test_writeARY(9'd127,16'b1010101010101010);

        test_writeARY(9'd128,16'b1100110011001100);
        test_writeARY(9'd129,16'b1100110011001100);
        test_writeARY(9'd130,16'b1100110011001100);
        test_writeARY(9'd131,16'b1100110011001100);
        test_writeARY(9'd132,16'b1100110011001100);
        test_writeARY(9'd133,16'b1100110011001100);
        test_writeARY(9'd134,16'b1100110011001100);
        test_writeARY(9'd135,16'b1100110011001100);
        test_writeARY(9'd136,16'b1100110011001100);
        test_writeARY(9'd137,16'b1100110011001100);
        test_writeARY(9'd138,16'b1100110011001100);
        test_writeARY(9'd139,16'b1100110011001100);
        test_writeARY(9'd140,16'b1100110011001100);
        test_writeARY(9'd141,16'b1100110011001100);
        test_writeARY(9'd142,16'b1100110011001100);
        test_writeARY(9'd143,16'b1100110011001100);
        test_writeARY(9'd144,16'b1100110011001100);
        test_writeARY(9'd145,16'b1100110011001100);
        test_writeARY(9'd146,16'b1100110011001100);
        test_writeARY(9'd147,16'b1100110011001100);
        test_writeARY(9'd148,16'b1100110011001100);
        test_writeARY(9'd149,16'b1100110011001100);
        test_writeARY(9'd150,16'b1100110011001100);
        test_writeARY(9'd151,16'b1100110011001100);
        test_writeARY(9'd152,16'b1100110011001100);
        test_writeARY(9'd153,16'b1100110011001100);
        test_writeARY(9'd154,16'b1100110011001100);
        test_writeARY(9'd155,16'b1100110011001100);
        test_writeARY(9'd156,16'b1100110011001100);
        test_writeARY(9'd157,16'b1100110011001100);
        test_writeARY(9'd158,16'b1100110011001100);
        test_writeARY(9'd159,16'b1100110011001100);
        test_writeARY(9'd160,16'b1100110011001100);
        test_writeARY(9'd161,16'b1100110011001100);
        test_writeARY(9'd162,16'b1100110011001100);
        test_writeARY(9'd163,16'b1100110011001100);
        test_writeARY(9'd164,16'b1100110011001100);
        test_writeARY(9'd165,16'b1100110011001100);
        test_writeARY(9'd166,16'b1100110011001100);
        test_writeARY(9'd167,16'b1100110011001100);
        test_writeARY(9'd168,16'b1100110011001100);
        test_writeARY(9'd169,16'b1100110011001100);
        test_writeARY(9'd170,16'b1100110011001100);
        test_writeARY(9'd171,16'b1100110011001100);
        test_writeARY(9'd172,16'b1100110011001100);
        test_writeARY(9'd173,16'b1100110011001100);
        test_writeARY(9'd174,16'b1100110011001100);
        test_writeARY(9'd175,16'b1100110011001100);
        test_writeARY(9'd176,16'b1100110011001100);
        test_writeARY(9'd177,16'b1100110011001100);
        test_writeARY(9'd178,16'b1100110011001100);
        test_writeARY(9'd179,16'b1100110011001100);
        test_writeARY(9'd180,16'b1100110011001100);
        test_writeARY(9'd181,16'b1100110011001100);
        test_writeARY(9'd182,16'b1100110011001100);
        test_writeARY(9'd183,16'b1100110011001100);
        test_writeARY(9'd184,16'b1100110011001100);
        test_writeARY(9'd185,16'b1100110011001100);
        test_writeARY(9'd186,16'b1100110011001100);
        test_writeARY(9'd187,16'b1100110011001100);
        test_writeARY(9'd188,16'b1100110011001100);
        test_writeARY(9'd189,16'b1100110011001100);
        test_writeARY(9'd190,16'b1100110011001100);
        test_writeARY(9'd191,16'b1100110011001100);
        test_writeARY(9'd192,16'b1100110011001100);
        test_writeARY(9'd193,16'b1100110011001100);
        test_writeARY(9'd194,16'b1100110011001100);
        test_writeARY(9'd195,16'b1100110011001100);
        test_writeARY(9'd196,16'b1100110011001100);
        test_writeARY(9'd197,16'b1100110011001100);
        test_writeARY(9'd198,16'b1100110011001100);
        test_writeARY(9'd199,16'b1100110011001100);
        test_writeARY(9'd200,16'b1100110011001100);
        test_writeARY(9'd201,16'b1100110011001100);
        test_writeARY(9'd202,16'b1100110011001100);
        test_writeARY(9'd203,16'b1100110011001100);
        test_writeARY(9'd204,16'b1100110011001100);
        test_writeARY(9'd205,16'b1100110011001100);
        test_writeARY(9'd206,16'b1100110011001100);
        test_writeARY(9'd207,16'b1100110011001100);
        test_writeARY(9'd208,16'b1100110011001100);
        test_writeARY(9'd209,16'b1100110011001100);
        test_writeARY(9'd210,16'b1100110011001100);
        test_writeARY(9'd211,16'b1100110011001100);
        test_writeARY(9'd212,16'b1100110011001100);
        test_writeARY(9'd213,16'b1100110011001100);
        test_writeARY(9'd214,16'b1100110011001100);
        test_writeARY(9'd215,16'b1100110011001100);
        test_writeARY(9'd216,16'b1100110011001100);
        test_writeARY(9'd217,16'b1100110011001100);
        test_writeARY(9'd218,16'b1100110011001100);
        test_writeARY(9'd219,16'b1100110011001100);
        test_writeARY(9'd220,16'b1100110011001100);
        test_writeARY(9'd221,16'b1100110011001100);
        test_writeARY(9'd222,16'b1100110011001100);
        test_writeARY(9'd223,16'b1100110011001100);
        test_writeARY(9'd224,16'b1100110011001100);
        test_writeARY(9'd225,16'b1100110011001100);
        test_writeARY(9'd226,16'b1100110011001100);
        test_writeARY(9'd227,16'b1100110011001100);
        test_writeARY(9'd228,16'b1100110011001100);
        test_writeARY(9'd229,16'b1100110011001100);
        test_writeARY(9'd230,16'b1100110011001100);
        test_writeARY(9'd231,16'b1100110011001100);
        test_writeARY(9'd232,16'b1100110011001100);
        test_writeARY(9'd233,16'b1100110011001100);
        test_writeARY(9'd234,16'b1100110011001100);
        test_writeARY(9'd235,16'b1100110011001100);
        test_writeARY(9'd236,16'b1100110011001100);
        test_writeARY(9'd237,16'b1100110011001100);
        test_writeARY(9'd238,16'b1100110011001100);
        test_writeARY(9'd239,16'b1100110011001100);
        test_writeARY(9'd240,16'b1100110011001100);
        test_writeARY(9'd241,16'b1100110011001100);
        test_writeARY(9'd242,16'b1100110011001100);
        test_writeARY(9'd243,16'b1100110011001100);
        test_writeARY(9'd244,16'b1100110011001100);
        test_writeARY(9'd245,16'b1100110011001100);
        test_writeARY(9'd246,16'b1100110011001100);
        test_writeARY(9'd247,16'b1100110011001100);
        test_writeARY(9'd248,16'b1100110011001100);
        test_writeARY(9'd249,16'b1100110011001100);
        test_writeARY(9'd250,16'b1100110011001100);
        test_writeARY(9'd251,16'b1100110011001100);
        test_writeARY(9'd252,16'b1100110011001100);
        test_writeARY(9'd253,16'b1100110011001100);
        test_writeARY(9'd254,16'b1100110011001100);
        test_writeARY(9'd255,16'b1100110011001100);

        test_writeARY(9'd256,16'b1111000011110000);
        test_writeARY(9'd257,16'b1111000011110000);
        test_writeARY(9'd258,16'b1111000011110000);
        test_writeARY(9'd259,16'b1111000011110000);
        test_writeARY(9'd260,16'b1111000011110000);
        test_writeARY(9'd261,16'b1111000011110000);
        test_writeARY(9'd262,16'b1111000011110000);
        test_writeARY(9'd263,16'b1111000011110000);
        test_writeARY(9'd264,16'b1111000011110000);
        test_writeARY(9'd265,16'b1111000011110000);
        test_writeARY(9'd266,16'b1111000011110000);
        test_writeARY(9'd267,16'b1111000011110000);
        test_writeARY(9'd268,16'b1111000011110000);
        test_writeARY(9'd269,16'b1111000011110000);
        test_writeARY(9'd270,16'b1111000011110000);
        test_writeARY(9'd271,16'b1111000011110000);
        test_writeARY(9'd272,16'b1111000011110000);
        test_writeARY(9'd273,16'b1111000011110000);
        test_writeARY(9'd274,16'b1111000011110000);
        test_writeARY(9'd275,16'b1111000011110000);
        test_writeARY(9'd276,16'b1111000011110000);
        test_writeARY(9'd277,16'b1111000011110000);
        test_writeARY(9'd278,16'b1111000011110000);
        test_writeARY(9'd279,16'b1111000011110000);
        test_writeARY(9'd280,16'b1111000011110000);
        test_writeARY(9'd281,16'b1111000011110000);
        test_writeARY(9'd282,16'b1111000011110000);
        test_writeARY(9'd283,16'b1111000011110000);
        test_writeARY(9'd284,16'b1111000011110000);
        test_writeARY(9'd285,16'b1111000011110000);
        test_writeARY(9'd286,16'b1111000011110000);
        test_writeARY(9'd287,16'b1111000011110000);
        test_writeARY(9'd288,16'b1111000011110000);
        test_writeARY(9'd289,16'b1111000011110000);
        test_writeARY(9'd290,16'b1111000011110000);
        test_writeARY(9'd291,16'b1111000011110000);
        test_writeARY(9'd292,16'b1111000011110000);
        test_writeARY(9'd293,16'b1111000011110000);
        test_writeARY(9'd294,16'b1111000011110000);
        test_writeARY(9'd295,16'b1111000011110000);
        test_writeARY(9'd296,16'b1111000011110000);
        test_writeARY(9'd297,16'b1111000011110000);
        test_writeARY(9'd298,16'b1111000011110000);
        test_writeARY(9'd299,16'b1111000011110000);
        test_writeARY(9'd300,16'b1111000011110000);
        test_writeARY(9'd301,16'b1111000011110000);
        test_writeARY(9'd302,16'b1111000011110000);
        test_writeARY(9'd303,16'b1111000011110000);
        test_writeARY(9'd304,16'b1111000011110000);
        test_writeARY(9'd305,16'b1111000011110000);
        test_writeARY(9'd306,16'b1111000011110000);
        test_writeARY(9'd307,16'b1111000011110000);
        test_writeARY(9'd308,16'b1111000011110000);
        test_writeARY(9'd309,16'b1111000011110000);
        test_writeARY(9'd310,16'b1111000011110000);
        test_writeARY(9'd311,16'b1111000011110000);
        test_writeARY(9'd312,16'b1111000011110000);
        test_writeARY(9'd313,16'b1111000011110000);
        test_writeARY(9'd314,16'b1111000011110000);
        test_writeARY(9'd315,16'b1111000011110000);
        test_writeARY(9'd316,16'b1111000011110000);
        test_writeARY(9'd317,16'b1111000011110000);
        test_writeARY(9'd318,16'b1111000011110000);
        test_writeARY(9'd319,16'b1111000011110000);
        test_writeARY(9'd320,16'b1111000011110000);
        test_writeARY(9'd321,16'b1111000011110000);
        test_writeARY(9'd322,16'b1111000011110000);
        test_writeARY(9'd323,16'b1111000011110000);
        test_writeARY(9'd324,16'b1111000011110000);
        test_writeARY(9'd325,16'b1111000011110000);
        test_writeARY(9'd326,16'b1111000011110000);
        test_writeARY(9'd327,16'b1111000011110000);
        test_writeARY(9'd328,16'b1111000011110000);
        test_writeARY(9'd329,16'b1111000011110000);
        test_writeARY(9'd330,16'b1111000011110000);
        test_writeARY(9'd331,16'b1111000011110000);
        test_writeARY(9'd332,16'b1111000011110000);
        test_writeARY(9'd333,16'b1111000011110000);
        test_writeARY(9'd334,16'b1111000011110000);
        test_writeARY(9'd335,16'b1111000011110000);
        test_writeARY(9'd336,16'b1111000011110000);
        test_writeARY(9'd337,16'b1111000011110000);
        test_writeARY(9'd338,16'b1111000011110000);
        test_writeARY(9'd339,16'b1111000011110000);
        test_writeARY(9'd340,16'b1111000011110000);
        test_writeARY(9'd341,16'b1111000011110000);
        test_writeARY(9'd342,16'b1111000011110000);
        test_writeARY(9'd343,16'b1111000011110000);
        test_writeARY(9'd344,16'b1111000011110000);
        test_writeARY(9'd345,16'b1111000011110000);
        test_writeARY(9'd346,16'b1111000011110000);
        test_writeARY(9'd347,16'b1111000011110000);
        test_writeARY(9'd348,16'b1111000011110000);
        test_writeARY(9'd349,16'b1111000011110000);
        test_writeARY(9'd350,16'b1111000011110000);
        test_writeARY(9'd351,16'b1111000011110000);
        test_writeARY(9'd352,16'b1111000011110000);
        test_writeARY(9'd353,16'b1111000011110000);
        test_writeARY(9'd354,16'b1111000011110000);
        test_writeARY(9'd355,16'b1111000011110000);
        test_writeARY(9'd356,16'b1111000011110000);
        test_writeARY(9'd357,16'b1111000011110000);
        test_writeARY(9'd358,16'b1111000011110000);
        test_writeARY(9'd359,16'b1111000011110000);
        test_writeARY(9'd360,16'b1111000011110000);
        test_writeARY(9'd361,16'b1111000011110000);
        test_writeARY(9'd362,16'b1111000011110000);
        test_writeARY(9'd363,16'b1111000011110000);
        test_writeARY(9'd364,16'b1111000011110000);
        test_writeARY(9'd365,16'b1111000011110000);
        test_writeARY(9'd366,16'b1111000011110000);
        test_writeARY(9'd367,16'b1111000011110000);
        test_writeARY(9'd368,16'b1111000011110000);
        test_writeARY(9'd369,16'b1111000011110000);
        test_writeARY(9'd370,16'b1111000011110000);
        test_writeARY(9'd371,16'b1111000011110000);
        test_writeARY(9'd372,16'b1111000011110000);
        test_writeARY(9'd373,16'b1111000011110000);
        test_writeARY(9'd374,16'b1111000011110000);
        test_writeARY(9'd375,16'b1111000011110000);
        test_writeARY(9'd376,16'b1111000011110000);
        test_writeARY(9'd377,16'b1111000011110000);
        test_writeARY(9'd378,16'b1111000011110000);
        test_writeARY(9'd379,16'b1111000011110000);
        test_writeARY(9'd380,16'b1111000011110000);
        test_writeARY(9'd381,16'b1111000011110000);
        test_writeARY(9'd382,16'b1111000011110000);
        test_writeARY(9'd383,16'b1111000011110000);

        test_writeARY(9'd384,16'b1111111100000000);
        test_writeARY(9'd385,16'b1111111100000000);
        test_writeARY(9'd386,16'b1111111100000000);
        test_writeARY(9'd387,16'b1111111100000000);
        test_writeARY(9'd388,16'b1111111100000000);
        test_writeARY(9'd389,16'b1111111100000000);
        test_writeARY(9'd390,16'b1111111100000000);
        test_writeARY(9'd391,16'b1111111100000000);
        test_writeARY(9'd392,16'b1111111100000000);
        test_writeARY(9'd393,16'b1111111100000000);
        test_writeARY(9'd394,16'b1111111100000000);
        test_writeARY(9'd395,16'b1111111100000000);
        test_writeARY(9'd396,16'b1111111100000000);
        test_writeARY(9'd397,16'b1111111100000000);
        test_writeARY(9'd398,16'b1111111100000000);
        test_writeARY(9'd399,16'b1111111100000000);
        test_writeARY(9'd400,16'b1111111100000000);
        test_writeARY(9'd401,16'b1111111100000000);
        test_writeARY(9'd402,16'b1111111100000000);
        test_writeARY(9'd403,16'b1111111100000000);
        test_writeARY(9'd404,16'b1111111100000000);
        test_writeARY(9'd405,16'b1111111100000000);
        test_writeARY(9'd406,16'b1111111100000000);
        test_writeARY(9'd407,16'b1111111100000000);
        test_writeARY(9'd408,16'b1111111100000000);
        test_writeARY(9'd409,16'b1111111100000000);
        test_writeARY(9'd410,16'b1111111100000000);
        test_writeARY(9'd411,16'b1111111100000000);
        test_writeARY(9'd412,16'b1111111100000000);
        test_writeARY(9'd413,16'b1111111100000000);
        test_writeARY(9'd414,16'b1111111100000000);
        test_writeARY(9'd415,16'b1111111100000000);
        test_writeARY(9'd416,16'b1111111100000000);
        test_writeARY(9'd417,16'b1111111100000000);
        test_writeARY(9'd418,16'b1111111100000000);
        test_writeARY(9'd419,16'b1111111100000000);
        test_writeARY(9'd420,16'b1111111100000000);
        test_writeARY(9'd421,16'b1111111100000000);
        test_writeARY(9'd422,16'b1111111100000000);
        test_writeARY(9'd423,16'b1111111100000000);
        test_writeARY(9'd424,16'b1111111100000000);
        test_writeARY(9'd425,16'b1111111100000000);
        test_writeARY(9'd426,16'b1111111100000000);
        test_writeARY(9'd427,16'b1111111100000000);
        test_writeARY(9'd428,16'b1111111100000000);
        test_writeARY(9'd429,16'b1111111100000000);
        test_writeARY(9'd430,16'b1111111100000000);
        test_writeARY(9'd431,16'b1111111100000000);
        test_writeARY(9'd432,16'b1111111100000000);
        test_writeARY(9'd433,16'b1111111100000000);
        test_writeARY(9'd434,16'b1111111100000000);
        test_writeARY(9'd435,16'b1111111100000000);
        test_writeARY(9'd436,16'b1111111100000000);
        test_writeARY(9'd437,16'b1111111100000000);
        test_writeARY(9'd438,16'b1111111100000000);
        test_writeARY(9'd439,16'b1111111100000000);
        test_writeARY(9'd440,16'b1111111100000000);
        test_writeARY(9'd441,16'b1111111100000000);
        test_writeARY(9'd442,16'b1111111100000000);
        test_writeARY(9'd443,16'b1111111100000000);
        test_writeARY(9'd444,16'b1111111100000000);
        test_writeARY(9'd445,16'b1111111100000000);
        test_writeARY(9'd446,16'b1111111100000000);
        test_writeARY(9'd447,16'b1111111100000000);
        test_writeARY(9'd448,16'b1111111100000000);
        test_writeARY(9'd449,16'b1111111100000000);
        test_writeARY(9'd450,16'b1111111100000000);
        test_writeARY(9'd451,16'b1111111100000000);
        test_writeARY(9'd452,16'b1111111100000000);
        test_writeARY(9'd453,16'b1111111100000000);
        test_writeARY(9'd454,16'b1111111100000000);
        test_writeARY(9'd455,16'b1111111100000000);
        test_writeARY(9'd456,16'b1111111100000000);
        test_writeARY(9'd457,16'b1111111100000000);
        test_writeARY(9'd458,16'b1111111100000000);
        test_writeARY(9'd459,16'b1111111100000000);
        test_writeARY(9'd460,16'b1111111100000000);
        test_writeARY(9'd461,16'b1111111100000000);
        test_writeARY(9'd462,16'b1111111100000000);
        test_writeARY(9'd463,16'b1111111100000000);
        test_writeARY(9'd464,16'b1111111100000000);
        test_writeARY(9'd465,16'b1111111100000000);
        test_writeARY(9'd466,16'b1111111100000000);
        test_writeARY(9'd467,16'b1111111100000000);
        test_writeARY(9'd468,16'b1111111100000000);
        test_writeARY(9'd469,16'b1111111100000000);
        test_writeARY(9'd470,16'b1111111100000000);
        test_writeARY(9'd471,16'b1111111100000000);
        test_writeARY(9'd472,16'b1111111100000000);
        test_writeARY(9'd473,16'b1111111100000000);
        test_writeARY(9'd474,16'b1111111100000000);
        test_writeARY(9'd475,16'b1111111100000000);
        test_writeARY(9'd476,16'b1111111100000000);
        test_writeARY(9'd477,16'b1111111100000000);
        test_writeARY(9'd478,16'b1111111100000000);
        test_writeARY(9'd479,16'b1111111100000000);
        test_writeARY(9'd480,16'b1111111100000000);
        test_writeARY(9'd481,16'b1111111100000000);
        test_writeARY(9'd482,16'b1111111100000000);
        test_writeARY(9'd483,16'b1111111100000000);
        test_writeARY(9'd484,16'b1111111100000000);
        test_writeARY(9'd485,16'b1111111100000000);
        test_writeARY(9'd486,16'b1111111100000000);
        test_writeARY(9'd487,16'b1111111100000000);
        test_writeARY(9'd488,16'b1111111100000000);
        test_writeARY(9'd489,16'b1111111100000000);
        test_writeARY(9'd490,16'b1111111100000000);
        test_writeARY(9'd491,16'b1111111100000000);
        test_writeARY(9'd492,16'b1111111100000000);
        test_writeARY(9'd493,16'b1111111100000000);
        test_writeARY(9'd494,16'b1111111100000000);
        test_writeARY(9'd495,16'b1111111100000000);
        test_writeARY(9'd496,16'b1111111100000000);
        test_writeARY(9'd497,16'b1111111100000000);
        test_writeARY(9'd498,16'b1111111100000000);
        test_writeARY(9'd499,16'b1111111100000000);
        test_writeARY(9'd500,16'b1111111100000000);
        test_writeARY(9'd501,16'b1111111100000000);
        test_writeARY(9'd502,16'b1111111100000000);
        test_writeARY(9'd503,16'b1111111100000000);
        test_writeARY(9'd504,16'b1111111100000000);
        test_writeARY(9'd505,16'b1111111100000000);
        test_writeARY(9'd506,16'b1111111100000000);
        test_writeARY(9'd507,16'b1111111100000000);
        test_writeARY(9'd508,16'b1111111100000000);
        test_writeARY(9'd509,16'b1111111100000000);
        test_writeARY(9'd510,16'b1111111100000000);
        test_writeARY(9'd511,16'b1111111100000000);
    //
    //calulation and read
        test_cal;
        test_read(5'd0,0);
        test_read(5'd1,0);
        test_read(5'd2,0);
        test_read(5'd3,0);
        test_read(5'd4,0);
        test_read(5'd5,0);
        test_read(5'd6,0);
        test_read(5'd7,0);
        test_read(5'd8,0);
        test_read(5'd9,0);
        test_read(5'd10,0);
        test_read(5'd11,0);
        test_read(5'd12,0);
        test_read(5'd13,0);
        test_read(5'd14,0);
        test_read(5'd15,0);
        # (CLK_PEROID*5);
    //
   // 
    // //test 2
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);



          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);

          
          test_writeBUF(5'd0,16'b1111111100000000);
          test_writeBUF(5'd1,16'b1111111100000000);
          test_writeBUF(5'd2,16'b0011001100110011);
          test_writeBUF(5'd3,16'b1111111111111111);
          test_writeBUF(5'd4,16'b1111111111111111);
          test_writeBUF(5'd5,16'b1111111111111111);
          test_writeBUF(5'd6,16'b1111111111111111);
          test_writeBUF(5'd7,16'b1111111111111111);
          test_writeBUF(5'd8,16'b1111111111111111);
          test_writeBUF(5'd9,16'b1111111111111111);
          test_writeBUF(5'd10,16'b1111111111111111);
          test_writeBUF(5'd11,16'b1111111111111111);
          test_writeBUF(5'd12,16'b1111111111111111);
          test_writeBUF(5'd13,16'b1111111111111111);
          test_writeBUF(5'd14,16'b1111111111111111);
          test_writeBUF(5'd15,16'b1111111111111111);
          test_writeBUF(5'd16,16'b1111111111111111);
          test_writeBUF(5'd17,16'b1111111111111111);
          test_writeBUF(5'd18,16'b1111111111111111);
          test_writeBUF(5'd19,16'b1111111111111111);
          test_writeBUF(5'd20,16'b1111111111111111);
          test_writeBUF(5'd21,16'b1111111111111111);
          test_writeBUF(5'd22,16'b1111111111111111);
          test_writeBUF(5'd23,16'b1111111111111111);
          test_writeBUF(5'd24,16'b1111111111111111);
          test_writeBUF(5'd25,16'b1111111111111111);
          test_writeBUF(5'd26,16'b1111111111111111);
          test_writeBUF(5'd27,16'b1111111111111111);
          test_writeBUF(5'd28,16'b1111111111111111);
          test_writeBUF(5'd29,16'b1111111111111111);
          test_writeBUF(5'd30,16'b1111111111111111);
          test_writeBUF(5'd31,16'b1111111111111111);

                  test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);


    // //
    // //test 3
    //       test_writeBUF(5'd0,16'b1111111100000000);
    //       test_writeBUF(5'd1,16'b1111111100000000);
    //       test_writeBUF(5'd2,16'b0011001100110011);
    //       test_writeBUF(5'd3,16'b1111111111111111);
    //       test_writeBUF(5'd4,16'b1111111111111111);
    //       test_writeBUF(5'd5,16'b1111111111111111);
    //       test_writeBUF(5'd6,16'b1111111111111111);
    //       test_writeBUF(5'd7,16'b1111111111111111);
    //       test_writeBUF(5'd8,16'b1111111111111111);
    //       test_writeBUF(5'd9,16'b1111111111111111);
    //       test_writeBUF(5'd10,16'b1111111111111111);
    //       test_writeBUF(5'd11,16'b1111111111111111);
    //       test_writeBUF(5'd12,16'b1111111111111111);
    //       test_writeBUF(5'd13,16'b1111111111111111);
    //       test_writeBUF(5'd14,16'b1111111111111111);
    //       test_writeBUF(5'd15,16'b1111111111111111);
    //       test_writeBUF(5'd16,16'b1111111111111111);
    //       test_writeBUF(5'd17,16'b1111111111111111);
    //       test_writeBUF(5'd18,16'b1111111111111111);
    //       test_writeBUF(5'd19,16'b1111111111111111);
    //       test_writeBUF(5'd20,16'b1111111111111111);
    //       test_writeBUF(5'd21,16'b1111111111111111);
    //       test_writeBUF(5'd22,16'b1111111111111111);
    //       test_writeBUF(5'd23,16'b1111111111111111);
    //       test_writeBUF(5'd24,16'b1111111111111111);
    //       test_writeBUF(5'd25,16'b1111111111111111);
    //       test_writeBUF(5'd26,16'b1111111111111111);
    //       test_writeBUF(5'd27,16'b1111111111111111);
    //       test_writeBUF(5'd28,16'b1111111111111111);
    //       test_writeBUF(5'd29,16'b1111111111111111);
    //       test_writeBUF(5'd30,16'b1111111111111111);
    //       test_writeBUF(5'd31,16'b1111111111111111);
    // //
    // //test 4
    //               test_cal;
    //       test_read(5'd0,0);
    //       test_read(5'd1,0);
    //       test_read(5'd2,0);
    //       test_read(5'd3,0);
    //       test_read(5'd4,0);
    //       test_read(5'd5,0);
    //       test_read(5'd6,0);
    //       test_read(5'd7,0);
    //       test_read(5'd8,0);
    //       test_read(5'd9,0);
    //       test_read(5'd10,0);
    //       test_read(5'd11,0);
    //       test_read(5'd12,0);
    //       test_read(5'd13,0);
    //       test_read(5'd14,0);
    //       test_read(5'd15,0);
    //       test_read(5'd16,0);
    //       test_read(5'd17,0);
    //       test_read(5'd18,0);
    //       test_read(5'd19,0);
    //       test_read(5'd20,0);
    //       test_read(5'd21,0);
    //       test_read(5'd22,0);
    //       test_read(5'd23,0);
    //       test_read(5'd24,0);
    //       test_read(5'd25,0);
    //       test_read(5'd26,0);
    //       test_read(5'd27,0);
    //       test_read(5'd28,0);
    //       test_read(5'd29,0);
    //       test_read(5'd30,0);
    //       test_read(5'd31,0);
    //       # (CLK_PEROID*5);

    //       test_writeBUF(5'd0,16'b1111111100000000);
    //       test_writeBUF(5'd1,16'b1111111100000000);
    //       test_writeBUF(5'd2,16'b0011001100110011);
    //       test_writeBUF(5'd3,16'b1111111111111111);
    //       test_writeBUF(5'd4,16'b1111111111111111);
    //       test_writeBUF(5'd5,16'b1111111111111111);
    //       test_writeBUF(5'd6,16'b1111111111111111);
    //       test_writeBUF(5'd7,16'b1111111111111111);
    //       test_writeBUF(5'd8,16'b1111111111111111);
    //       test_writeBUF(5'd9,16'b1111111111111111);
    //       test_writeBUF(5'd10,16'b1111111111111111);
    //       test_writeBUF(5'd11,16'b1111111111111111);
    //       test_writeBUF(5'd12,16'b1111111111111111);
    //       test_writeBUF(5'd13,16'b1111111111111111);
    //       test_writeBUF(5'd14,16'b1111111111111111);
    //       test_writeBUF(5'd15,16'b1111111111111111);
    //       test_writeBUF(5'd16,16'b1111111111111111);
    //       test_writeBUF(5'd17,16'b1111111111111111);
    //       test_writeBUF(5'd18,16'b1111111111111111);
    //       test_writeBUF(5'd19,16'b1111111111111111);
    //       test_writeBUF(5'd20,16'b1111111111111111);
    //       test_writeBUF(5'd21,16'b1111111111111111);
    //       test_writeBUF(5'd22,16'b1111111111111111);
    //       test_writeBUF(5'd23,16'b1111111111111111);
    //       test_writeBUF(5'd24,16'b1111111111111111);
    //       test_writeBUF(5'd25,16'b1111111111111111);
    //       test_writeBUF(5'd26,16'b1111111111111111);
    //       test_writeBUF(5'd27,16'b1111111111111111);
    //       test_writeBUF(5'd28,16'b1111111111111111);
    //       test_writeBUF(5'd29,16'b1111111111111111);
    //       test_writeBUF(5'd30,16'b1111111111111111);
    //       test_writeBUF(5'd31,16'b1111111111111111);

    //       test_cal;
    //       test_read(5'd0,0);
    //       test_read(5'd1,0);
    //       test_read(5'd2,0);
    //       test_read(5'd3,0);
    //       test_read(5'd4,0);
    //       test_read(5'd5,0);
    //       test_read(5'd6,0);
    //       test_read(5'd7,0);
    //       test_read(5'd8,0);
    //       test_read(5'd9,0);
    //       test_read(5'd10,0);
    //       test_read(5'd11,0);
    //       test_read(5'd12,0);
    //       test_read(5'd13,0);
    //       test_read(5'd14,0);
    //       test_read(5'd15,0);
    //       test_read(5'd16,0);
    //       test_read(5'd17,0);
    //       test_read(5'd18,0);
    //       test_read(5'd19,0);
    //       test_read(5'd20,0);
    //       test_read(5'd21,0);
    //       test_read(5'd22,0);
    //       test_read(5'd23,0);
    //       test_read(5'd24,0);
    //       test_read(5'd25,0);
    //       test_read(5'd26,0);
    //       test_read(5'd27,0);
    //       test_read(5'd28,0);
    //       test_read(5'd29,0);
    //       test_read(5'd30,0);
    //       test_read(5'd31,0);
    //       # (CLK_PEROID*5);
    // //
    // //test 5
    //       test_writeBUF(5'd0,16'b1111111100000000);
    //       test_writeBUF(5'd1,16'b1000110000001110);
    //       test_writeBUF(5'd2,16'b0011001100110000);
    //       test_writeBUF(5'd3,16'b1110111101000001);
    //       test_writeBUF(5'd4,16'b1000101110011001);
    //       test_writeBUF(5'd5,16'b1111111111111111);
    //       test_writeBUF(5'd6,16'b1100111100000011);
    //       test_writeBUF(5'd7,16'b1111111111111111);
    //       test_writeBUF(5'd8,16'b1101111100001101);
    //       test_writeBUF(5'd9,16'b1111111111111111);
    //       test_writeBUF(5'd10,16'b1111111111111111);
    //       test_writeBUF(5'd11,16'b1111111111111111);
    //       test_writeBUF(5'd12,16'b1111111011111111);
    //       test_writeBUF(5'd13,16'b1001011111100011);
    //       test_writeBUF(5'd14,16'b1111111000111110);
    //       test_writeBUF(5'd15,16'b1111111111111111);
    //       test_writeBUF(5'd16,16'b1111111111111111);
    //       test_writeBUF(5'd17,16'b1111000011101111);
    //       test_writeBUF(5'd19,16'b1111111111111111);
    //       test_writeBUF(5'd20,16'b1111111111111111);
    //       test_writeBUF(5'd21,16'b1111111111111111);
    //       test_writeBUF(5'd22,16'b1111111111110010);
    //       test_writeBUF(5'd23,16'b1111011010000011);
    //       test_writeBUF(5'd25,16'b1111111110011111);
    //       test_writeBUF(5'd26,16'b1100111111110001);
    //       test_writeBUF(5'd27,16'b1111111111111001);
    //       test_writeBUF(5'd28,16'b1110011111000000);
    //       test_writeBUF(5'd29,16'b1111111110000111);
    //       test_writeBUF(5'd30,16'b1110011111111001);
    //       test_writeBUF(5'd31,16'b1110010001111111);

    //               test_cal;
    //       test_read(5'd0,0);
    //       test_read(5'd1,0);
    //       test_read(5'd2,0);
    //       test_read(5'd3,0);
    //       test_read(5'd4,0);
    //       test_read(5'd5,0);
    //       test_read(5'd6,0);
    //       test_read(5'd7,0);
    //       test_read(5'd8,0);
    //       test_read(5'd9,0);
    //       test_read(5'd10,0);
    //       test_read(5'd11,0);
    //       test_read(5'd12,0);
    //       test_read(5'd13,0);
    //       test_read(5'd14,0);
    //       test_read(5'd15,0);
    //       test_read(5'd16,0);
    //       test_read(5'd17,0);
    //       test_read(5'd18,0);
    //       test_read(5'd19,0);
    //       test_read(5'd20,0);
    //       test_read(5'd21,0);
    //       test_read(5'd22,0);
    //       test_read(5'd23,0);
    //       test_read(5'd24,0);
    //       test_read(5'd25,0);
    //       test_read(5'd26,0);
    //       test_read(5'd27,0);
    //       test_read(5'd28,0);
    //       test_read(5'd29,0);
    //       test_read(5'd30,0);
    //       test_read(5'd31,0);
    //       # (CLK_PEROID*5);
    // //
    // //test 6
    //       test_writeBUF(5'd0,16'b1111111100000000);
    //       test_writeBUF(5'd1,16'b1111111100000000);
    //       test_writeBUF(5'd2,16'b0011001100110011);
    //       test_writeBUF(5'd3,16'b1111111001000011);
    //       test_writeBUF(5'd4,16'b1110000111110011);
    //       test_writeBUF(5'd5,16'b1111111111111111);
    //       test_writeBUF(5'd6,16'b1111111111000011);
    //       test_writeBUF(5'd7,16'b0011100111100111);
    //       test_writeBUF(5'd8,16'b1111001111100011);
    //       test_writeBUF(5'd9,16'b11111100001111111);
    //       test_writeBUF(5'd10,16'b1111111111111001);
    //       test_writeBUF(5'd11,16'b1111110001111111);
    //       test_writeBUF(5'd12,16'b1111001111110110);
    //       test_writeBUF(5'd13,16'b1111111111111111);
    //       test_writeBUF(5'd14,16'b1111111000011111);
    //       test_writeBUF(5'd15,16'b1001111111100111);
    //       test_writeBUF(5'd16,16'b0111110011111111);
    //       test_writeBUF(5'd17,16'b1001111111100001);
    //       test_writeBUF(5'd18,16'b1111001110011111);
    //       test_writeBUF(5'd19,16'b1111111111111111);
    //       test_writeBUF(5'd20,16'b1111111000011111);
    //       test_writeBUF(5'd21,16'b1110011111100111);
    //       test_writeBUF(5'd22,16'b1111111111111111);
    //       test_writeBUF(5'd23,16'b1110011111111111);
    //       test_writeBUF(5'd24,16'b1111111111111111);
    //       test_writeBUF(5'd25,16'b1111111000111111);
    //       test_writeBUF(5'd26,16'b1111111111111111);
    //       test_writeBUF(5'd27,16'b1100001111111111);
    //       test_writeBUF(5'd28,16'b1111111111100001);
    //       test_writeBUF(5'd29,16'b1001111001110011);
    //       test_writeBUF(5'd30,16'b1111001111111111);
    //       test_writeBUF(5'd31,16'b1100001111100111);

    //               test_cal;
    //       test_read(5'd0,0);
    //       test_read(5'd1,0);
    //       test_read(5'd2,0);
    //       test_read(5'd3,0);
    //       test_read(5'd4,0);
    //       test_read(5'd5,0);
    //       test_read(5'd6,0);
    //       test_read(5'd7,0);
    //       test_read(5'd8,0);
    //       test_read(5'd9,0);
    //       test_read(5'd10,0);
    //       test_read(5'd11,0);
    //       test_read(5'd12,0);
    //       test_read(5'd13,0);
    //       test_read(5'd14,0);
    //       test_read(5'd15,0);
    //       test_read(5'd16,0);
    //       test_read(5'd17,0);
    //       test_read(5'd18,0);
    //       test_read(5'd19,0);
    //       test_read(5'd20,0);
    //       test_read(5'd21,0);
    //       test_read(5'd22,0);
    //       test_read(5'd23,0);
    //       test_read(5'd24,0);
    //       test_read(5'd25,0);
    //       test_read(5'd26,0);
    //       test_read(5'd27,0);
    //       test_read(5'd28,0);
    //       test_read(5'd29,0);
    //       test_read(5'd30,0);
    //       test_read(5'd31,0);
    
   
    //test 7
        test_writeBUF(5'd0,16'b0000000000000000);
        test_writeBUF(5'd1,16'b0000000000000000);
        test_writeBUF(5'd2,16'b0000000000000000);
        test_writeBUF(5'd3,16'b0000000000000000);
        test_writeBUF(5'd4,16'b0000000000000000);
        test_writeBUF(5'd5,16'b0000000000000000);
        test_writeBUF(5'd6,16'b0000000000000000);
        test_writeBUF(5'd7,16'b0000000000000000);
        test_writeBUF(5'd8,16'b0000000000000000);
        test_writeBUF(5'd9,16'b0000000000000000);
        test_writeBUF(5'd10,16'b0000000000000000);
        test_writeBUF(5'd11,16'b0000000000000000);
        test_writeBUF(5'd12,16'b0000000000000000);
        test_writeBUF(5'd13,16'b0000000000000000);
        test_writeBUF(5'd14,16'b0000000000000000);
        test_writeBUF(5'd15,16'b0000000000000000);
        test_writeBUF(5'd16,16'b0000000000000000);
        test_writeBUF(5'd17,16'b0000000000000000);
        test_writeBUF(5'd18,16'b0000000000000000);
        test_writeBUF(5'd19,16'b0000000000000000);
        test_writeBUF(5'd20,16'b0000000000000000);
        test_writeBUF(5'd21,16'b0000000000000000);
        test_writeBUF(5'd22,16'b0000000000000000);
        test_writeBUF(5'd23,16'b0000000000000000);
        test_writeBUF(5'd24,16'b0000000000000000);
        test_writeBUF(5'd25,16'b0000000000000000);
        test_writeBUF(5'd26,16'b0000000000000000);
        test_writeBUF(5'd27,16'b0000000000000000);
        test_writeBUF(5'd28,16'b0000000000000000);
        test_writeBUF(5'd29,16'b0000000000000000);
        test_writeBUF(5'd30,16'b0000000000000000);
        test_writeBUF(5'd31,16'b0000000000000000);

          test_cal;
          test_read(5'd0,0);
          test_read(5'd1,0);
          test_read(5'd2,0);
          test_read(5'd3,0);
          test_read(5'd4,0);
          test_read(5'd5,0);
          test_read(5'd6,0);
          test_read(5'd7,0);
          test_read(5'd8,0);
          test_read(5'd9,0);
          test_read(5'd10,0);
          test_read(5'd11,0);
          test_read(5'd12,0);
          test_read(5'd13,0);
          test_read(5'd14,0);
          test_read(5'd15,0);
          # (CLK_PEROID*5);
    //
    //
    $finish(10);
        
    end


endmodule