* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
***************************************************************************************** 
* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for HSPICE only)  
*****************************************************************************************
*
* Release version    : 1.11
*
* Release date       : 4/30/2015
*
* Simulation tool    : Synopsys Star-HSPICE version 2006.09
*
*
*   MOSFET Varactor  :
*
*        *----------------------------------------------------------------------* 
*        |                      MOSFET varactor subckt                          |
*        |======================================================================| 
*        |   NMOS in NWELL 1.8V      | pvar18_ckt_rf                            | 
*        |======================================================================| 
*        |   NMOS in NWELL 3.3V      | pvar33_ckt_rf                            | 
*        *----------------------------------------------------------------------*
*
*   
*   Junction Diode Varactor  :
*
*        *----------------------------------------------------------------------* 
*        | Junction Diode type       |               1.8V | 3.3V                |
*        |======================================================================| 
*        |          N+/PWELL         |     pvardio18_rf   |    pvardio33_rf     |
*        *----------------------------------------------------------------------*
* 
*        *----------------------------------------------------------------------* 
*        | Junction Diode subckt     |               1.8V | 3.3V                |
*        |======================================================================| 
*        |          N+/PWELL         |   pvardio18_ckt_rf | pvardio33_ckt_rf    |
*        *----------------------------------------------------------------------*
*
*            
***************************
* 0.18um 1.8V MOS Varactor*
***************************
* 1=port1, 2=port2
* Area=wr*lr*nf
.subckt pvar18_ckt_rf 1 2 lr=l wr=w nf=finger mr=1 mismod_var=1
* 1.8v mos varactor scalable model parameters
.param
**mismatch parameter
+ac0_pvar18_rf     =  0          
+bc0_pvar18_rf     =  3.04e-9    
+cc0_pvar18_rf     =  0  
+geo_var_rf        = 'ac0_pvar18_rf/(wr*(lr+2.6e-14/lr)*nf*mr)+bc0_pvar18_rf/sqrt(wr*(lr+2.6e-14/lr)*nf*mr)+cc0_pvar18_rf'         
+dcgg_pvar18mis_rf = 'mismod_var*sigma_mis_var_rf*geo_var_rf' 
**subckt parameter              
+rsub1_rf     = 'max((-629.32*log(nf)+4000), 1e-3)' 
+csub1_rf     = 'max((0.0348*nf+0.1652)*1e-15, 1e-18)'
+cox1_rf      = 'max(((0.004*(lr*1e6)+0.0081)*(wr*1e6)*nf+(0.032*(lr*1e6)+0.0638))*1e-15, 1e-18)'
+rsub2_rf     = 'max((303.64*(lr*1e6)+254.47)*pwr((wr*1e6)*nf,(-0.3054*(lr*1e6)+0.0147)), 1e-3)'
+csub2_rf     = 'max((((0.8728*(lr*1e6)-0.528)*(wr*1e6)+(-3.1644*(lr*1e6)+4.2208))*nf+((-1.7148*(lr*1e6)+4.3055)*(wr*1e6)+(0.6456*(lr*1e6)+1.4517)))*1e-15, 1e-18)'
+cox2_rf      = 'max((((0.126*(lr*1e6)+0.0168)*(wr*1e6)+(0.896*(lr*1e6)+0.828))*nf+((-0.0204*(lr*1e6)+1.4385)*(wr*1e6)+(-0.163*(lr*1e6)+1.0508)))*1e-15, 1e-18)'
+djnw_area_rf = '(wr*1e6+2*0.12)*(lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*1e-12'
+djnw_pj_rf   = '(wr*1e6+2*0.12+lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*2*1e-6'
+cgg_a2       = 'a_a2*((8.28*(wr*1e6)*(lr*1e6)*nf+0.4638*(wr*1e6)*nf+0.7149*(lr*1e6)*nf+0.202*(wr*1e6)-0.1569*(lr*1e6)))'
+cgg_a1       = 'a_a1*((1.647*(wr*1e6)*(lr*1e6)*nf+0.4773*(wr*1e6)*nf+0.5422*(lr*1e6)*nf+0.04776*(wr*1e6)+0.01854*(lr*1e6)))'
+cgg_x0       = '-0.4315*pwr((wr*1e6),-0.07108)*(1-2.758*(lr*1e6)+1.902*(lr*1e6)*(lr*1e6))*pwr(nf+552.3,0.07095*pwr((wr*1e6),0.01743)*pwr((lr*1e6),-1.0097))'
+a_a1	      = '1.0704*exp(-0.0385*(lr*1e6))'
+a_a2	      = '0.0361*log(lr*1e6)+0.9651'
+rs_rf        = 'max((((((-7.562e-01*(lr*1e6)+1.839e+00)*(wr*1e6)*(wr*1e6)+(6.514e+00*(lr*1e6)-2.316e+01)*(wr*1e6)+(-3.931e+01*(lr*1e6)+1.370e+02))*pwr(nf,((4.100e-03*(lr*1e6)-4.300e-03)*(wr*1e6)*(wr*1e6)+(-4.590e-02*(lr*1e6)+4.900e-02)*(wr*1e6)+(1.446e-01*(lr*1e6)-1.153e+00))))))*(1+drs_pvar18_rf), 1e-6)'
**gate current parameter
+tox    = '1.2518e-08+dtox_pvar18_rf' 
+gcie   = 2.449260179                 gcarc = 4.97112503779554                 gcevgc = 1.28405488039671
+gcetc  = 2425.31845182089            gcete = 0.305811750223937                igg_tc = 0.00896             
gg  22 2 current='((v(22,2)*pwr(abs(v(22,2)),gcie)*(gcarc*wr*(lr+2.6e-14/lr)*nf*exp(gcevgc*v(22,2)-gcetc*pwr(tox,gcete))))*1)*(1+igg_tc*(temper-25))' m=mr
* equivalent circuit
ls    11 22  10p       m=mr    
rs    1  11  r = 'max((((rs_rf*(1+0.04/(v(22,2)*v(22,2)+(0.0004*(wr*1e6)*(wr*1e6)+0.0137*(wr*1e6)+0.4708)*(0.0004*(wr*1e6)*(wr*1e6)+0.0137*(wr*1e6)+0.4708))))*(1+2.266e-03*(temper-25)-3.309e-06*(temper-25)*(temper-25)))), 1e-6)' m=mr          
cgg   22  2  c='max((cgg_a2+(cgg_a1-cgg_a2)/(1+exp((v(22,2)-cgg_x0)/((-0.0347*v(22,2)*v(22,2)*v(22,2)*v(22,2)+0.00857*v(22,2)*v(22,2)*v(22,2)+0.131*v(22,2)*v(22,2)-0.0389*v(22,2)+0.19)*(0.00143*(temper-25)+1)))))*(1+dcgg_pvar18_rf)*1e-15, 1e-15)' m=mr
cox1  1  10  cox1_rf   m=mr 
rsub1 10  0  rsub1_rf  m=mr 
csub1 10  0  csub1_rf  m=mr 
cox2  2  20  cox2_rf   m=mr     
rsub2 20  0  rsub2_rf  m=mr 
csub2 20  0  csub2_rf  m=mr 
djnw  0   2
+nwdio_rf
+area  = djnw_area_rf
+pj    = djnw_pj_rf   
+m     = mr      
.model  nwdio_rf  d  level = 3
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+dcap    = 2               area    = 9.6e-009        pj      = 4e-004          tref    = 25
**************************************************************
*               DC PARAMETERS
**************************************************************
+is      = 2.3733e-006     jsw     = 2.9142e-014                vb      = 15              ibv     = 104
+ikr     = 104170          n       = 1.085                      rs      = 8.4602e-009
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+cj      = 0               cjp     = 0               pb      = 0.41624         php     = 0.81575
+fcs     = 0               mj      = 0.26295         mjsw    = 0.377           fc      = 0
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+tlev    = 1               tlevc   = 1               trs     = 0.0004       xti     = 3
+cta     = 0.0017608       ctp     = 0.0012659       tpb     = 0.00155      tphp    = 0.0022128
+eg      = 1.16
*
.ends pvar18_ckt_rf
*
*************************************
* 0.18um 3.3V MOS Varactor
*************************************
* 1=port1, 2=port2
* Area=wr*lr*nf
.subckt pvar33_ckt_rf 1 2 lr=l wr=w nf=finger mr=1  mismod_var=1
.param
*+Ar         = 'lr*wr*nf'    
*+Ls_rf      = 'max(((-2.32720800*lr*1e6+3.84952400)*pwr(wr*1e6*nf,(-0.02020000*lr*1e6-0.96951500)))*1E-9, 1E-15)'
+Rsub1_rf   = 'max((-157.33*log(nf)+1000), 1E-3)'
+Csub1_rf   = 'max(((0.058000*lr*1e6+0.131000)*nf+(1.152200*lr*1e6+0.263900))*1E-15, 1E-18)'
+Cox1_rf    = 'max((((-0.02130818*lr*1e6+0.02299185)*wr*1e6+(0.19167958*lr*1e6-0.03172040))*nf+(-0.01930408*lr*1e6+0.02256428)*wr*1e6+(0.03578980*lr*1e6-0.12376429))*1E-15, 1E-18)'
+Rsub2_rf   = 'max(((0.17509600*lr*1e6+0.13622500)*wr*1e6+(-3.13181000*lr*1e6-5.98751100))*nf+(-0.36204000*lr*1e6-16.93326600)*wr*1e6+(-5.25510200*lr*1e6+ 419.97183700), 1E-3)'
+Csub2_rf   = 'max((((-0.05913800*lr*1e6+3.56503100)*wr*1e6+(2.06525200*lr*1e6+0.32525500))*pwr(nf,((0.02163000*lr*1e6-0.05084700)*wr*1e6+(-0.18202800*lr*1e6+0.69376000))))*1E-15, 1E-18)'
+Cox2_rf    = 'max((((0.03803200*lr*1e6+0.07406700)*wr*1e6+(1.19708000*lr*1e6+0.60749200))*nf+(0.10622800*lr*1e6+1.37163800)*wr*1e6+(-0.25722800*lr*1e6+1.02081900))*1E-15, 1E-18)'
+Djnw_AREA_rf = '(wr*1e6+2*0.12)*(lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*1e-12'
+Djnw_PJ_rf   = '(wr*1e6+2*0.12+lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*2*1e-6'
+Rs_A = '(((2.18219600*lr*1e6-1.31073200)*wr*1e6*wr*1e6+(-36.30831000*lr*1e6+23.46962700)*wr*1e6+(106.27523200*lr*1e6-24.91322400))*pwr(nf,((-0.02877400*lr*1e6+0.02830400)*wr*1e6*wr*1e6+(0.40768000*lr*1e6-0.40029000)*wr*1e6+(-1.23126600*lr*1e6+0.17806600))))'
+Rs_B = '((-0.56984200*lr*1e6+0.59987600)*wr*1e6*wr*1e6+(8.46208200*lr*1e6-9.01834500)*wr*1e6+(-27.19727400*lr*1e6+30.22506800))'
+Rs_D = '((-0.05474200*lr*1e6+0.05283200)*wr*1e6*wr*1e6+(0.80293400*lr*1e6-0.77210600)*wr*1e6+(-2.13486200*lr*1e6+2.90342700))'
+Rs_E = '((-0.02549600*lr*1e6+0.03906600)*wr*1e6*wr*1e6+(0.48609400*lr*1e6-0.70076400)*wr*1e6+(-2.59254400*lr*1e6+3.40643400))'
+Cgg_A1     = 'a_a1*((4.924416E+00*lr*1e6+3.885705E-01)*a_a1w*wr*1e6*nf+(5.756613E-02*lr*1e6+3.680246E-01))'
+Cgg_A2     = 'a_a2*((1.490944E+00*lr*1e6+4.324138E-01)*a_a2w*wr*1e6*nf+(-9.410417E-02*lr*1e6+3.779284E-01))'
+Cgg_x0     = '(-(-2.510018E-02*lr*1e6+2.329891E-01)*pwr(wr*1e6*nf,(2.091532E-02*lr*1e6-2.966834E-02)))'
+Cgg_dx     = '(-(3.454607E-02*lr*1e6+3.079878E-01)*pwr(wr*1e6*nf,(-1.125777E-02*lr*1e6+2.882598E-03)))'
+a_a1	= '1.0147*pwr(wr*1e6,-0.0211)'
+a_a2	= '1.0+0.0157*log(nf)'
+a_a1w	= 1
+a_a2w	= 1
*** mismatch paramters	
+lrr='lr*1e6' wrr='wr*1e6'     
+area = 'lrr*wrr*nf'        
+geo_var_rf = 'ac0_pvar33_rf/sqrt(area*mr)+bc0_pvar33_rf'	
+dcgg_pvar33mis_rf = 'mismod_var*sigma_mis_var_rf*geo_var_rf'
* equivalent circuit
Ls    11 22  10p    m=mr
Rs    1  11  R= 'max(((Rs_A*(1+0.1*Rs_E*V(22,2)+0.1*Rs_B/(V(22,2)*V(22,2)+Rs_D*Rs_D)))*(1+2.266E-03*(temper-25)-3.309E-06*(temper-25)*(temper-25)))*(1+DRS_PVAR33_RF),1E-6)' m=mr
Rsub1 10  0  Rsub1_rf m=mr
Csub1 10  0  Csub1_rf m=mr
Cox1  1  10  Cox1_rf  m=mr
Rsub2 20  0  Rsub2_rf m=mr
Csub2 20  0  Csub2_rf m=mr
Djnw  0 2
+ nwdio_rf
+ AREA  = Djnw_AREA_rf
+ PJ    = Djnw_PJ_rf
+ m     = mr
Cox2  2  20  Cox2_rf m=mr
Cgg   22  2  C='max(((Cgg_A2+(Cgg_A1-Cgg_A2)/(1+EXP((V(22,2)-Cgg_x0)/(Cgg_dx*(0.00143*(temper-25)+1))))))*(1+dcgg_pvar33mis_rf)*(1+DCGG_PVAR33_RF)*1e-15, 1e-15)' m=mr
*.model nwdio_rf d
*+LEVEL    = 3                   JS       = 1.42E-06            JSW      = 1.00E-15            
*+N        = 1.0128              RS       = 2.44E-08            IK       = 1.1E+04            
*+IKR      = 1.04E+05            BV       = 15.0                IBV      = 104.2               
*+TRS      = 9.47E-04            EG       = 1.16                TREF     = 25.0                
*+XTI      = 3.0                 CJ       = 0           MJ       = 0.317               
*+PB       = 0.494               CJSW     = 0               MJSW     = 0.383               
*+PHP      = 0.9                 CTA      = 0.002               CTP      = 0.00121                 
*+TPB      = 0.00253             TPHP     = 0.00217             TLEV     = 1
*+TLEVC    = 1    FC       = 0                   FCS      = 0                
.model  nwdio_rf  d  level = 3
**************************************************************
*               GENERAL PARAMETERS
**************************************************************
+dcap    = 2               area    = 9.6e-009        pj      = 4e-004          tref    = 25
**************************************************************
*               DC PARAMETERS
**************************************************************
+is      = 2.3733e-006     jsw     = 2.9142e-014     vb      = 15              ibv     = 104
+ikr     = 104170          n       = 1.085           rs      = 8.4602e-009
**************************************************************
*               CAPACITANCE PARAMETERS
**************************************************************
+cj      = 0        cjp     = 0     pb      = 0.41624         php     = 0.81575
+fcs     = 0        mj      = 0.26295         mjsw    = 0.377           fc      = 0
**************************************************************
*               NOISE PARAMETERS
**************************************************************
**************************************************************
*               TEMPERATURE PARAMETERS
**************************************************************
+tlev    = 1               tlevc   = 1               trs     = 0.0004       xti     = 3
+cta     = 0.0017608       ctp     = 0.0012659       tpb     = 0.00155      tphp    = 0.0022128
+eg      = 1.16
.ends pvar33_ckt_rf
*
****************************
* 0.18um 1.8V P+/NW Varactor
****************************
* 1=port1, 2=port2
* Area=wr*lr*nf
.subckt pvardio18_ckt_rf 1 2 lr=l wr=w nf=finger
* P+/NW junction varactor scalable model parameters
.param
+Ar        = 'lr*wr*nf'
+Pj        = '(lr+wr)*2*nf'
+Ls_rf     = '(0.07947+(1.7134E-05*Ar*1E12)-(3.865E-09*Ar*Ar*1E24))*1E-9'
+Rs_rf     = '0.23268+(3.334E+03/(Ar*1E12))+(8.9147E+04/(Ar*Ar*1E24))'
+Rsub1_rf  = '1E+5'
+Csub1_rf  = '1*1E-15'
+Cox1_rf   = '1*1E-15'
+Rsub2_rf  = '1940-(1.6342*Ar*1E12)+(4.2816E-04*Ar*Ar*1E24)'
+Csub2_rf  = '(2.75025+(2.787E-03*Ar*1E12)+(1.3682E-06*Ar*Ar*1E24))*1E-15'
+Cox2_rf   = '(27.96263+(0.53519*Ar*1E12)-(9.0589E-05*Ar*Ar*1E24))*1E-15'
Ls    1 11    LS_rf        
Rs    11 22   Rs_rf    
Cox1  1 10  Cox1_rf  
Csub1 10 0 Csub1_rf
Rsub1 10 0 Rsub1_rf        
Cox2  2 20  Cox2_rf  
Csub2 20 0 Csub2_rf
Rsub2 20 0 Rsub2_rf
Diode 22 2 pvardio18_rf AREA=Ar PJ=Pj
* P+/Nwell varactor Model
.MODEL pvardio18_rf D
+LEVEL   = 3            CJ   = 1.1495E-3          MJ    = 0.37316    
+TREF    = 25           PB   = 0.76958            CTA   = 0.000876
+TPB     = 0.00153      FC   = 0                  FCS   = 0              
+EG      = 1.16         TLEV = 1                  TLEVC = 1   
+JS       = 1.1913E-07            JSW      = 1e-15            
+N        = 0.98812              RS       = 0           IK     = 4.2216e+06            
+IKR      = 2000000            BV       = 12                IBV    = 2000            
+TRS      = 1.78E-03           XTI      = 3.0                 
.ends pvardio18_ckt_rf
*
****************************
* 0.18um 3.3V P+/NW Varactor
****************************
* 1=port1, 2=port2
* Area=wr*lr*nf
.subckt pvardio33_ckt_rf 1 2 lr=l wr=w nf=finger
* P+/NW junction varactor scalable model parameters
.param
+Ar        = 'lr*wr*nf'
+Pj        = '(lr+wr)*2*nf'
+Ls_rf     = '(0.08203+(1.3302E-05*Ar*1E12)-(1.844E-09*Ar*Ar*1E24))*1E-9' 
+Rs_rf     = '0.25902+(3.3475E+03/(Ar*1E12))+(1.0295E+05/(Ar*Ar*1E24))'
+Rsub1_rf  = '1E+5'
+Csub1_rf  = '1*1E-15'
+Cox1_rf   = '1*1E-15'
+Rsub2_rf  = '1.869E+03-(1.49373*Ar*1E12)+(3.7877E-04*Ar*Ar*1E24)'
+Csub2_rf  = '(3.81691-(1.5322E-03*Ar*1E12)+(4.0789E-06*Ar*Ar*1E24))*1E-15'
+Cox2_rf   = '(64.90675+(0.37036*Ar*1E12)+(1.0985E-06*Ar*Ar*1E24))*1E-15'
Ls    1 11    LS_rf        
Rs    11 22   Rs_rf    
Cox1  1 10  Cox1_rf  
Csub1 10 0 Csub1_rf
Rsub1 10 0 Rsub1_rf        
Cox2  2 20  Cox2_rf  
Csub2 20 0 Csub2_rf
Rsub2 20 0 Rsub2_rf
Diode 22 2 pvardio33_rf AREA=Ar PJ=Pj
* P+/Nwell varactor Model
.MODEL pvardio33_rf D
+LEVEL   = 3            CJ   = 1.1455E-3          MJ    = 0.3793    
+TREF    = 25           PB   = 0.792              CTA   = 0.000897
+TPB     = 0.00166      FC   = 0                  FCS   = 0
+EG      = 1.16         TLEV = 1                  TLEVC = 1
+JS       = 1.3141E-07            JSW      = 1E-15             
+N        = 0.99195             RS       = 0            IK       = 4.5171E+06            
+IKR      = 2000000            BV       = 12                IBV      = 2000              
+TRS      = 1.24E-03           XTI      = 3.0                 
.ends pvardio33_ckt_rf
