* 
* No part of this file can be released without the consent of SMIC.
*
************************************************************************************************************
* smic 0.18um mixed signal 1p6m 1.8v/3.3v spice model(for HSPICE only) *
************************************************************************************************************
*
* Release version    : 1.11
*
* Release date       : 18/03/2015
*
* Simulation tool    : Synopsys Star-HSPICE version C-2009.09
*
*  Inductor   :
* *  *------------------------*---------------------------------------------------------*
*    |  Turn, Radius & Width  |  T=2~7.5 step 0.5,W=3~15um,R=1.7071*W+11.878~120um       |
* *  *------------------------*---------------------------------------------------------*
*    |        Model Name      |              diff_ind_rf_psub                           |
* *  *------------------------*---------------------------------------------------------*
.subckt diff_ind_rf_psub PLUS MINUS PSUB R=6e-05 w=8e-06 n=3
.param radius_='0.00833333*(R/1e-06-0)' w_='0.0666667*(w/1e-06-0)'
.param T54='(1-abs(sgn(n-(2.5))))'
.param T55='(min(sgn(radius_-(0.416958))+1,1))'
.param T56='(min(sgn(w_-(0.6004))+1,1))'
.param T57='(min(sgn(w_-(0.5996))+1,1))'
.param T58='(min(sgn(radius_-(0.416375))+1,1))'
.param T59='(min(sgn(radius_-(0.708625))+1,1))'
.param T60='(min(sgn(radius_-(0.708042))+1,1))'
.param T61='(1-abs(sgn(n-(2))))'
.param T62='(1-abs(sgn(n-(3.5))))'
.param T63='(1-abs(sgn(n-(3))))'
.param T64='(1-abs(sgn(n-(4.5))))'
.param T65='(1-abs(sgn(n-(4))))'
.param T66='(1-abs(sgn(n-(5.5))))'
.param T67='(1-abs(sgn(n-(5))))'
.param T68='(1-abs(sgn(n-(6.5))))'
.param T69='(1-abs(sgn(n-(6))))'
.param T70='(1-abs(sgn(n-(7.5))))'
.param T71='(1-abs(sgn(n-(7))))'
.param S0='T54*(1-T55)*(1-T56)'
.param noS0='(1-S0)'
.param S1='T54*T57*(1-T55)*noS0'
.param noS1='(1-S1)*noS0'
.param S2='T54*(1-T56)*T58*(1-T59)*noS1'
.param noS2='(1-S2)*noS1'
.param S3='T54*T58*T57*(1-T59)*noS2'
.param noS3='(1-S3)*noS2'
.param S4='T54*(1-T56)*T60*noS3'
.param noS4='(1-S4)*noS3'
.param S5='T54*T60*T57*noS4'
.param noS5='(1-S5)*noS4'
.param S6='T61*(1-T55)*(1-T56)*noS5'
.param noS6='(1-S6)*noS5'
.param S7='T61*T57*(1-T55)*noS6'
.param noS7='(1-S7)*noS6'
.param S8='T61*(1-T56)*T58*(1-T59)*noS7'
.param noS8='(1-S8)*noS7'
.param S9='T61*T58*T57*(1-T59)*noS8'
.param noS9='(1-S9)*noS8'
.param S10='T61*(1-T56)*T60*noS9'
.param noS10='(1-S10)*noS9'
.param S11='T61*T60*T57*noS10'
.param noS11='(1-S11)*noS10'
.param S12='T62*(1-T55)*noS11'
.param noS12='(1-S12)*noS11'
.param S13='T62*T58*(1-T59)*noS12'
.param noS13='(1-S13)*noS12'
.param S14='T62*T60*noS13'
.param noS14='(1-S14)*noS13'
.param S15='T63*(1-T55)*(1-T56)*noS14'
.param noS15='(1-S15)*noS14'
.param S16='T63*T57*(1-T55)*noS15'
.param noS16='(1-S16)*noS15'
.param S17='T63*(1-T56)*T58*(1-T59)*noS16'
.param noS17='(1-S17)*noS16'
.param S18='T63*T58*T57*(1-T59)*noS17'
.param noS18='(1-S18)*noS17'
.param S19='T63*(1-T56)*T60*noS18'
.param noS19='(1-S19)*noS18'
.param S20='T63*T60*T57*noS19'
.param noS20='(1-S20)*noS19'
.param S21='T64*(1-T55)*noS20'
.param noS21='(1-S21)*noS20'
.param S22='T64*T58*(1-T59)*noS21'
.param noS22='(1-S22)*noS21'
.param S23='T64*T60*noS22'
.param noS23='(1-S23)*noS22'
.param S24='T65*(1-T55)*noS23'
.param noS24='(1-S24)*noS23'
.param S25='T65*T58*(1-T59)*noS24'
.param noS25='(1-S25)*noS24'
.param S26='T65*T60*noS25'
.param noS26='(1-S26)*noS25'
.param S27='T66*(1-T55)*noS26'
.param noS27='(1-S27)*noS26'
.param S28='T66*T58*(1-T59)*noS27'
.param noS28='(1-S28)*noS27'
.param S29='T66*T60*noS28'
.param noS29='(1-S29)*noS28'
.param S30='T67*(1-T55)*noS29'
.param noS30='(1-S30)*noS29'
.param S31='T67*T58*(1-T59)*noS30'
.param noS31='(1-S31)*noS30'
.param S32='T67*T60*noS31'
.param noS32='(1-S32)*noS31'
.param S33='T68*(1-T55)*noS32'
.param noS33='(1-S33)*noS32'
.param S34='T68*T58*(1-T59)*noS33'
.param noS34='(1-S34)*noS33'
.param S35='T68*T60*noS34'
.param noS35='(1-S35)*noS34'
.param S36='T69*(1-T55)*noS35'
.param noS36='(1-S36)*noS35'
.param S37='T69*T58*(1-T59)*noS36'
.param noS37='(1-S37)*noS36'
.param S38='T69*T60*noS37'
.param noS38='(1-S38)*noS37'
.param S39='T70*(1-T55)*noS38'
.param noS39='(1-S39)*noS38'
.param S40='T70*T58*(1-T59)*noS39'
.param noS40='(1-S40)*noS39'
.param S41='T70*T60*noS40'
.param noS41='(1-S41)*noS40'
.param S42='T71*(1-T55)*noS41'
.param noS42='(1-S42)*noS41'
.param S43='T71*T58*(1-T59)*noS42'
.param noS43='(1-S43)*noS42'
.param S44='T71*T60*noS43'
.param noS44='(1-S44)*noS43'
.param V0_part1='(-2.077232e+00)*S0+(-1.912155e-01)*S1+1.437538e+00*S2+(-4.361856e-01)*S3+(-8.423784e-02)*S4+2.408252e+00*S5+0.000000e+00*S6+1.795240e+00*S7+0.000000e+00*S8+(-2.267216e+00)*S9'
.param V0_part2='V0_part1+2.774136e+00*S10+(-1.326970e+01)*S11+(-8.428740e-02)*S12+3.639081e+00*S13+(-5.468273e+00)*S14+2.507956e-01*S15+3.788856e+00*S16+1.829262e+00*S17+7.366488e+00*S18+3.764977e-01*S19'
.param V0_part3='V0_part2+1.352043e+01*S20+8.016475e-01*S21+3.505367e+00*S22+1.822467e-01*S23+3.289699e+00*S24+(-1.492827e+00)*S25+7.128410e+00*S26+5.791254e+00*S27+5.157686e+00*S28+1.890551e+00*S29'
.param V0_part4='V0_part3+5.178105e+00*S30+5.858419e+00*S31+6.121661e+00*S32+(-2.379717e-01)*S33+4.827852e+00*S34+8.463019e+00*S35+8.201781e+00*S36+(-1.229384e+01)*S37+(-1.330177e-01)*S38+1.082419e+01*S39'
.param V0='V0_part4+8.073163e-02*S40+1.666474e-01*S41+7.996847e+00*S42+2.747680e+00*S43+(-3.605014e-01)*S44'
.param V1_part1='3.557242e+01*S0+2.050977e+01*S1+2.734904e+01*S2+3.833343e+01*S3+3.533548e+01*S4+3.323144e+01*S5+0.000000e+00*S6+9.444727e+00*S7+0.000000e+00*S8+1.534621e+01*S9'
.param V1_part2='V1_part1+6.259691e+00*S10+3.107095e+01*S11+5.590457e+01*S12+5.033975e+01*S13+6.962645e+01*S14+2.725020e+01*S15+3.170059e+01*S16+3.407847e+01*S17+2.562174e+01*S18+3.188559e+01*S19'
.param V1_part3='V1_part2+2.070987e+01*S20+7.608561e+01*S21+7.105378e+01*S22+9.278282e+01*S23+5.497211e+01*S24+8.562493e+01*S25+5.332130e+01*S26+1.026700e+02*S27+1.055221e+02*S28+1.252967e+02*S29'
.param V1_part4='V1_part3+8.383528e+01*S30+7.753407e+01*S31+7.699003e+01*S32+1.476813e+02*S33+1.394557e+02*S34+1.210593e+02*S35+1.087822e+02*S36+1.578081e+02*S37+1.326773e+02*S38+1.628431e+02*S39'
.param V1='V1_part4+1.894469e+02*S40+1.660640e+02*S41+1.426656e+02*S42+1.548591e+02*S43+1.632845e+02*S44'
.param V2_part1='4.563072e+00*S0+1.097208e+01*S1+(-1.044569e+00)*S2+(-3.340752e+00)*S3+(-2.118428e+00)*S4+(-1.489286e-01)*S5+0.000000e+00*S6+(-2.216679e+00)*S7+0.000000e+00*S8+4.494775e+00*S9'
.param V2_part2='V2_part1+5.104752e+00*S10+(-7.657718e-01)*S11+2.340432e+00*S12+(-8.645128e+00)*S13+1.096578e+01*S14+8.572361e+00*S15+4.604986e+00*S16+(-9.334558e+00)*S17+(-8.505680e+00)*S18+(-2.030521e+00)*S19'
.param V2_part3='V2_part2+(-1.399522e+01)*S20+1.780164e+01*S21+1.715537e+01*S22+1.784834e+00*S23+(-6.666806e+00)*S24+9.078933e+00*S25+(-1.081230e+01)*S26+8.731836e+00*S27+(-1.147156e+00)*S28+1.474750e+01*S29'
.param V2_part4='V2_part3+(-1.984505e+00)*S30+1.449485e+01*S31+1.172236e+01*S32+7.207681e+01*S33+1.989913e+00*S34+1.629093e+01*S35+6.861830e+00*S36+7.913137e+01*S37+3.278323e+01*S38+2.641047e+01*S39'
.param V2='V2_part4+6.760988e+01*S40+1.530341e+01*S41+1.858122e+01*S42+(-1.783179e+00)*S43+5.641521e+01*S44'
.param V3_part1='2.089292e+01*S0+(-2.873297e-01)*S1+(-1.085887e+00)*S2+(-6.562453e-01)*S3+(-1.337298e+00)*S4+(-1.679749e+00)*S5+(-9.165562e-01)*S6+2.036357e-01*S7+(-1.299786e+00)*S8+(-2.189496e+00)*S9'
.param V3_part2='V3_part1+4.563259e-01*S10+(-1.263891e+00)*S11+(-3.144424e+00)*S12+(-2.958244e+00)*S13+(-3.586912e+00)*S14+3.319352e+01*S15+1.273820e+01*S16+(-1.651952e+00)*S17+(-7.716882e-01)*S18+(-3.787381e-02)*S19'
.param V3_part3='V3_part2+(-1.808344e+00)*S20+4.559898e+00*S21+9.309684e+01*S22+(-1.784679e+01)*S23+(-1.060994e+00)*S24+(-3.487110e+00)*S25+3.389168e+01*S26+(-2.359234e+00)*S27+(-3.145759e+00)*S28+(-4.347432e+01)*S29'
.param V3_part4='V3_part3+(-1.158532e+00)*S30+(-3.397456e+00)*S31+(-6.049750e+00)*S32+(-1.508346e+00)*S33+4.023971e+03*S34+9.845788e+03*S35+(-1.615391e+00)*S36+(-4.943028e+00)*S37+(-6.684534e+01)*S38+(-1.461311e+00)*S39'
.param V3='V3_part4+1.264906e+02*S40+(-1.019337e+01)*S41+(-1.478845e+00)*S42+(-3.398639e+00)*S43+(-5.769078e+01)*S44'
.param V4_part1='(-6.804268e+01)*S0+1.294997e+00*S1+3.235921e+00*S2+2.017533e+00*S3+(-8.738561e-02)*S4+2.695749e+00*S5+6.790303e+00*S6+3.580765e-01*S7+(-8.349746e-01)*S8+9.546499e-01*S9'
.param V4_part2='V4_part1+(-6.626049e+00)*S10+5.085588e-01*S11+(-3.006775e+00)*S12+1.097419e+01*S13+1.353787e+00*S14+(-9.395303e+01)*S15+(-2.240036e+01)*S16+5.140542e+00*S17+2.415598e+00*S18+(-1.427146e+00)*S19'
.param V4_part3='V4_part2+3.108826e+00*S20+6.105686e+01*S21+2.517184e+02*S22+4.093075e+01*S23+1.046255e+01*S24+1.881680e+00*S25+1.734021e+02*S26+4.536347e-02*S27+3.128887e+00*S28+1.208827e+02*S29'
.param V4_part4='V4_part3+1.418900e+01*S30+8.829016e+00*S31+9.081465e+00*S32+2.358608e+01*S33+3.431269e+02*S34+1.964552e+02*S35+3.583221e-02*S36+2.323869e+01*S37+1.826386e+02*S38+3.154871e+00*S39'
.param V4='V4_part4+2.775570e+02*S40+1.949475e+01*S41+2.425214e+01*S42+3.816000e+00*S43+1.598358e+02*S44'
.param V5_part1='2.670730e+01*S0+4.806980e-01*S1+6.397334e-01*S2+6.422539e-01*S3+2.960482e+00*S4+1.120314e+00*S5+2.623207e-01*S6+1.157126e+00*S7+3.217394e+00*S8+7.995361e+00*S9'
.param V5_part2='V5_part1+7.766722e+00*S10+3.021387e+00*S11+4.864918e+00*S12+8.876290e-01*S13+4.813169e+00*S14+2.654107e+01*S15+4.459583e+01*S16+7.560944e-01*S17+7.547997e-01*S18+3.298603e+00*S19'
.param V5_part3='V5_part2+1.216922e+00*S20+(-8.771613e-01)*S21+(-3.426022e+01)*S22+1.573278e+00*S23+5.377527e-01*S24+3.830209e+00*S25+(-2.469923e+01)*S26+4.513043e+00*S27+3.740415e+00*S28+(-8.705960e-01)*S29'
.param V5_part4='V5_part3+6.834938e-01*S30+1.264536e+00*S31+1.859279e+00*S32+1.022618e+00*S33+(-8.230544e+02)*S34+(-1.975270e+03)*S35+4.114718e+00*S36+1.443920e+00*S37+(-3.099414e+00)*S38+3.985495e+00*S39'
.param V5='V5_part4+(-3.075017e+01)*S40+3.117689e+00*S41+1.051173e+00*S42+4.606575e+00*S43+(-1.204461e+00)*S44'
.param V6_part1='(-1.524699e-01)*S0+(-3.824031e-02)*S1+(-9.056454e-02)*S2+(-5.359134e-02)*S3+5.811417e-02*S4+(-1.069326e-01)*S5+(-2.339148e-02)*S6+3.165152e-03*S7+1.153322e-01*S8+(-8.829582e-03)*S9'
.param V6_part2='V6_part1+6.409554e-01*S10+7.745771e-02*S11+8.945718e-02*S12+(-2.253696e-01)*S13+(-1.842834e-01)*S14+(-1.445640e-01)*S15+5.949245e-02*S16+(-1.079534e-01)*S17+(-6.259764e-02)*S18+3.816822e-01*S19'
.param V6_part3='V6_part2+(-1.859525e-01)*S20+(-2.159284e-01)*S21+(-7.961430e+00)*S22+(-7.059345e-01)*S23+(-7.230197e-02)*S24+1.044219e-02*S25+(-6.570348e+00)*S26+2.024240e-02*S27+(-6.433422e-02)*S28+(-1.564415e+00)*S29'
.param V6_part4='V6_part3+(-1.045914e-01)*S30+(-4.431617e-01)*S31+(-7.452344e-01)*S32+(-1.506952e-01)*S33+(-9.794701e+00)*S34+(-2.411411e+01)*S35+1.801043e-04*S36+(-3.198724e-01)*S37+(-2.311028e+00)*S38+1.149333e-02*S39'
.param V6='V6_part4+4.980484e+00*S40+(-6.168724e-01)*S41+(-1.427875e-01)*S42+(-2.240520e-01)*S43+(-2.680388e+00)*S44'
.param V7_part1='8.312163e+00*S0+1.664494e+00*S1+2.044237e+00*S2+1.821156e+00*S3+1.933292e+00*S4+2.107675e+00*S5+1.116328e+00*S6+9.148044e-01*S7+1.015364e+00*S8+1.432942e+00*S9'
.param V7_part2='V7_part1+9.748282e-01*S10+1.069684e+00*S11+2.861165e+00*S12+3.929784e+00*S13+3.966923e+00*S14+1.061769e+01*S15+1.105903e+01*S16+2.630284e+00*S17+2.314208e+00*S18+2.331131e+00*S19'
.param V7_part3='V7_part2+2.692687e+00*S20+6.221335e+00*S21+3.968788e+01*S22+7.175245e+00*S23+3.943831e+00*S24+4.069612e+00*S25+1.624512e+01*S26+6.469744e+00*S27+7.380151e+00*S28+1.092768e+01*S29'
.param V7_part4='V7_part3+5.944773e+00*S30+6.665670e+00*S31+7.339017e+00*S32+1.000727e+01*S33+1.883149e+01*S34+2.353763e+01*S35+7.286906e+00*S36+9.454819e+00*S37+1.277818e+01*S38+1.126121e+01*S39'
.param V7='V7_part4+1.562682e+01*S40+1.548850e+01*S41+1.101653e+01*S42+1.093467e+01*S43+1.607835e+01*S44'
.param V8_part1='7.171267e-02*S0+(-2.700319e-03)*S1+(-9.836715e-02)*S2+(-2.341447e-02)*S3+(-5.057312e-01)*S4+(-1.617940e-01)*S5+(-2.358715e-02)*S6+(-4.177379e-02)*S7+(-2.298918e-01)*S8+(-8.645159e-02)*S9'
.param V8_part2='V8_part1+(-7.005024e-01)*S10+(-2.032071e-01)*S11+(-2.398407e-01)*S12+(-5.005919e-02)*S13+(-1.033338e+00)*S14+(-3.820925e-02)*S15+(-4.364340e-01)*S16+(-1.026122e-01)*S17+(-2.984918e-02)*S18+(-8.793217e-01)*S19'
.param V8_part3='V8_part2+(-1.672065e-01)*S20+1.993605e-01*S21+7.375369e+00*S22+(-6.756903e-01)*S23+4.959381e-02*S24+(-6.477498e-01)*S25+8.210229e+00*S26+6.891022e-02*S27+(-5.524374e-01)*S28+(-3.133667e-02)*S29'
.param V8_part4='V8_part3+3.126237e-01*S30+5.185575e-01*S31+2.232677e-01*S32+1.185233e+00*S33+3.849484e+01*S34+7.821247e+01*S35+2.151026e-01*S36+4.522650e-02*S37+6.973959e-01*S38+1.050005e+00*S39'
.param V8='V8_part4+(-1.301139e+00)*S40+(-1.612990e+00)*S41+1.370614e+00*S42+(-1.613009e-01)*S43+1.364726e+00*S44'
.param V9_part1='(-1.108868e+00)*S0+1.937720e+01*S1+(-4.016642e+00)*S2+(-4.171624e+00)*S3+(-9.123212e+00)*S4+(-6.630886e-01)*S5+(-1.963667e+00)*S6+(-9.868120e-01)*S7+(-2.036483e+00)*S8+(-8.926941e-01)*S9'
.param V9_part2='V9_part1+(-3.292705e+00)*S10+(-2.474757e+00)*S11+(-1.972513e+00)*S12+(-6.470472e+00)*S13+(-1.051368e+01)*S14+(-1.273683e+00)*S15+(-5.474439e-01)*S16+(-2.260604e+00)*S17+(-2.465540e+00)*S18+(-1.106341e+01)*S19'
.param V9_part3='V9_part2+(-2.329596e+00)*S20+(-2.784100e+00)*S21+(-4.833631e+00)*S22+(-6.257438e+00)*S23+(-3.567333e+00)*S24+(-6.711411e+00)*S25+(-6.779276e+00)*S26+(-2.319907e+00)*S27+(-1.092587e+01)*S28+(-7.392413e+00)*S29'
.param V9_part4='V9_part3+(-4.587418e+00)*S30+7.643392e+01*S31+1.207810e+02*S32+(-2.962641e+00)*S33+(-4.701424e+00)*S34+(-8.569964e+00)*S35+(-2.904024e+00)*S36+(-7.106669e+00)*S37+(-7.691075e+00)*S38+(-2.792103e+00)*S39'
.param V9='V9_part4+(-4.660892e+00)*S40+(-3.127231e+00)*S41+(-3.121526e+00)*S42+(-1.342032e+01)*S43+(-9.311526e+00)*S44'
.param V10_part1='5.656080e+00*S0+(-4.855655e+01)*S1+(-1.570155e+00)*S2+7.528411e-01*S3+1.645855e+01*S4+1.731350e-02*S5+2.674136e+00*S6+3.971595e+00*S7+5.498524e+00*S8+2.170044e+00*S9'
.param V10_part2='V10_part1+4.737464e+00*S10+4.164944e+00*S11+1.552400e+01*S12+3.178688e+00*S13+1.836627e+01*S14+6.548824e+00*S15+2.881736e+00*S16+(-6.206129e-01)*S17+1.262509e+00*S18+1.791824e+01*S19'
.param V10_part3='V10_part2+4.616901e-01*S20+9.651876e+00*S21+8.682899e+00*S22+5.308378e+00*S23+(-1.098583e+00)*S24+2.355536e+01*S25+7.247187e+00*S26+3.183088e+01*S27+5.227062e+01*S28+8.234547e+00*S29'
.param V10_part4='V10_part3+1.154608e+00*S30+(-1.835007e+02)*S31+(-1.862437e+02)*S32+2.717128e+00*S33+1.059059e+01*S34+1.108150e+01*S35+3.800113e+01*S36+5.100264e+00*S37+9.007333e+00*S38+6.419647e+01*S39'
.param V10='V10_part4+1.292635e+01*S40+(-1.816441e+01)*S41+1.701279e+00*S42+6.402371e+01*S43+1.025922e+01*S44'
.param V11_part1='7.656152e-01*S0+5.854812e+01*S1+1.011923e+01*S2+1.147589e+01*S3+2.068111e+00*S4+7.701474e+00*S5+2.028362e+00*S6+8.652880e-01*S7+9.579124e-01*S8+9.810576e-01*S9'
.param V11_part2='V11_part1+1.424924e+00*S10+1.535643e+00*S11+1.024258e+00*S12+6.817512e+00*S13+3.116477e+00*S14+8.587734e-01*S15+1.044488e+00*S16+6.960763e+00*S17+1.022385e+01*S18+2.637866e+00*S19'
.param V11_part3='V11_part2+9.702942e+00*S20+2.343391e+00*S21+3.025859e+00*S22+6.194200e+00*S23+6.651792e+00*S24+2.011748e+00*S25+3.755931e+00*S26+1.627551e+00*S27+2.730302e+00*S28+5.922338e+00*S29'
.param V11_part4='V11_part3+7.758870e+00*S30+4.263483e+01*S31+5.274095e+01*S32+8.040276e+00*S33+4.267744e+00*S34+5.868279e+00*S35+1.770436e+00*S36+9.304537e+00*S37+5.955718e+00*S38+2.377971e+00*S39'
.param V11='V11_part4+4.669207e+00*S40+2.814132e+01*S41+8.887051e+00*S42+3.929251e+00*S43+7.540718e+00*S44'
.param V12_part1='(-6.144087e-02)*S0+3.126460e-01*S1+4.381914e-01*S2+4.749843e-01*S3+(-3.040343e-01)*S4+3.608020e-01*S5+(-1.506915e-02)*S6+(-3.111807e-02)*S7+(-5.026159e-02)*S8+(-8.101660e-02)*S9'
.param V12_part2='V12_part1+(-1.493173e-01)*S10+(-1.995526e-01)*S11+(-1.156528e-01)*S12+1.090188e-01*S13+(-8.478783e-01)*S14+(-9.145272e-02)*S15+(-1.038399e-01)*S16+3.826183e-01*S17+3.963377e-01*S18+(-5.173121e-01)*S19'
.param V12_part3='V12_part2+3.813797e-01*S20+3.086638e-01*S21+2.421625e-01*S22+(-2.645982e-01)*S23+4.608906e-04*S24+(-4.340751e-01)*S25+2.855886e-02*S26+(-2.447840e-01)*S27+(-8.835723e-01)*S28+(-3.735981e-01)*S29'
.param V12_part4='V12_part3+(-1.028076e-02)*S30+1.507902e+00*S31+(-1.768212e-01)*S32+1.472347e-02*S33+8.001949e-02*S34+(-3.460489e-01)*S35+(-2.574551e-01)*S36+(-1.829545e-01)*S37+(-4.484235e-01)*S38+(-3.233534e-01)*S39'
.param V12='V12_part4+3.779985e-01*S40+(-1.207860e+00)*S41+1.925166e-02*S42+(-7.391321e-01)*S43+(-5.136353e-01)*S44'
.param V13_part1='3.581687e+00*S0+1.168421e+01*S1+3.594940e+00*S2+3.166783e+00*S3+4.671392e+00*S4+3.448859e+00*S5+1.980472e+00*S6+2.082678e+00*S7+2.383872e+00*S8+2.174833e+00*S9'
.param V13_part2='V13_part1+2.689174e+00*S10+2.548837e+00*S11+6.479128e+00*S12+6.607428e+00*S13+8.831708e+00*S14+4.572610e+00*S15+4.206038e+00*S16+4.351441e+00*S17+4.113732e+00*S18+6.274883e+00*S19'
.param V13_part3='V13_part2+4.531736e+00*S20+9.300381e+00*S21+1.049713e+01*S22+1.154993e+01*S23+6.983847e+00*S24+9.249230e+00*S25+8.956790e+00*S26+1.474387e+01*S27+1.745361e+01*S28+1.656215e+01*S29'
.param V13_part4='V13_part3+1.049535e+01*S30+5.117770e+01*S31+5.914462e+01*S32+1.746175e+01*S33+2.008315e+01*S34+2.232411e+01*S35+1.661232e+01*S36+1.650070e+01*S37+1.863905e+01*S38+2.588933e+01*S39'
.param V13='V13_part4+2.539609e+01*S40+2.747518e+01*S41+1.928611e+01*S42+2.455730e+01*S43+2.443533e+01*S44'
.param V14_part1='(-9.574332e-02)*S0+(-2.593114e-01)*S1+(-8.009068e-01)*S2+(-5.118057e-01)*S3+(-6.329866e-01)*S4+(-6.504260e-01)*S5+(-1.417353e-01)*S6+(-4.642940e-02)*S7+(-2.090779e-01)*S8+(-8.490650e-02)*S9'
.param V14_part2='V14_part1+(-4.657057e-01)*S10+(-1.595815e-01)*S11+9.386906e-02*S12+(-1.142969e+00)*S13+(-1.296274e+00)*S14+(-9.707723e-02)*S15+2.675117e-02*S16+(-8.576154e-01)*S17+(-5.173813e-01)*S18+(-7.696210e-01)*S19'
.param V14_part3='V14_part2+(-8.617898e-01)*S20+(-2.197990e-01)*S21+(-1.110977e+00)*S22+(-2.487675e+00)*S23+(-2.881161e-01)*S24+(-3.415344e-01)*S25+(-1.969979e+00)*S26+1.146449e+00*S27+4.251655e-01*S28+(-3.033971e+00)*S29'
.param V14_part4='V14_part3+(-6.811822e-02)*S30+(-7.390063e+00)*S31+(-1.256175e+01)*S32+9.221517e-01*S33+(-7.948418e-01)*S34+(-3.235248e+00)*S35+1.485201e+00*S36+(-9.596572e-01)*S37+(-3.119450e+00)*S38+4.057782e+00*S39'
.param V14='V14_part4+(-4.136599e-01)*S40+(-2.609107e+00)*S41+1.268894e+00*S42+9.478426e-01*S43+(-3.333939e+00)*S44'
.param V15_part1='(-2.257574e-01)*S0+(-3.449851e-01)*S1+2.519909e-01*S2+(-1.896722e-01)*S3+(-3.705675e-01)*S4+(-8.610797e-02)*S5+1.790918e-01*S6+5.467518e-01*S7+(-9.239621e-02)*S8+3.687930e-01*S9'
.param V15_part2='V15_part1+(-2.854786e-01)*S10+2.378390e-01*S11+(-1.750818e-01)*S12+2.660884e-01*S13+3.015592e+00*S14+(-2.466618e-01)*S15+(-5.456384e-01)*S16+(-4.584471e-03)*S17+(-1.149429e-01)*S18+(-3.739737e-01)*S19'
.param V15_part3='V15_part2+1.242477e-01*S20+3.803790e-01*S21+(-9.348190e-01)*S22+7.221089e-01*S23+(-1.317906e-01)*S24+8.486879e-01*S25+1.431141e-01*S26+3.833578e-02*S27+1.300365e+00*S28+(-2.450142e+01)*S29'
.param V15_part4='V15_part3+(-2.920200e-02)*S30+(-9.431010e-02)*S31+6.520289e-03*S32+2.180114e-01*S33+(-2.237242e+00)*S34+2.120297e+01*S35+6.099120e-03*S36+(-8.530409e-01)*S37+1.156473e-01*S38+2.634775e-01*S39'
.param V15='V15_part4+(-1.517581e+00)*S40+4.719027e+02*S41+7.451821e-02*S42+2.861881e+03*S43+1.000000e+04*S44'
.param V16_part1='5.266506e-01*S0+4.455534e-01*S1+8.151304e-01*S2+1.163855e+00*S3+3.031947e+00*S4+1.164366e+00*S5+6.420254e+00*S6+1.430499e+00*S7+1.761566e+00*S8+7.846322e-02*S9'
.param V16_part2='V16_part1+7.811655e-01*S10+9.455030e-01*S11+4.318080e+00*S12+2.686712e+00*S13+(-9.066390e-01)*S14+7.337639e-01*S15+7.639468e-01*S16+1.615053e+00*S17+1.250180e+00*S18+1.366557e+00*S19'
.param V16_part3='V16_part2+9.155497e-01*S20+6.571884e-01*S21+1.665209e+00*S22+4.511807e+00*S23+6.152482e+00*S24+1.610282e+00*S25+2.548710e-01*S26+6.246488e+00*S27+3.831750e+00*S28+3.609637e+01*S29'
.param V16_part4='V16_part3+6.549667e+00*S30+9.010835e-01*S31+5.023910e-01*S32+7.220144e+00*S33+3.571777e+00*S34+2.007683e+03*S35+7.572911e+00*S36+8.423792e+00*S37+1.299803e+02*S38+7.692991e+00*S39'
.param V16='V16_part4+2.672145e+00*S40+8.772362e+02*S41+7.886482e+00*S42+4.112866e+02*S43+1.000000e+04*S44'
.param V17_part1='(-2.264018e+00)*S0+(-6.784873e-01)*S1+(-3.024832e-01)*S2+1.392523e-01*S3+(-2.081939e-01)*S4+2.311639e-02*S5+2.844550e-01*S6+5.164612e-02*S7+(-2.571795e-02)*S8+(-2.712553e-01)*S9'
.param V17_part2='V17_part1+(-7.486064e-03)*S10+(-8.486067e-02)*S11+1.352241e-01*S12+(-1.904060e-01)*S13+(-1.436275e+00)*S14+(-2.338170e+00)*S15+(-1.122653e+00)*S16+(-1.059100e-02)*S17+1.662101e-01*S18+2.801829e-01*S19'
.param V17_part3='V17_part2+1.288395e-01*S20+(-5.341458e-01)*S21+(-1.984732e+00)*S22+4.377694e-01*S23+1.182300e+00*S24+(-8.247064e-02)*S25+(-1.296564e+00)*S26+1.102034e+00*S27+9.306564e-02*S28+2.921668e+01*S29'
.param V17_part4='V17_part3+1.180714e+00*S30+(-3.068496e+00)*S31+(-3.069520e+00)*S32+1.234002e+00*S33+6.589686e+00*S34+2.262904e+02*S35+1.162374e+00*S36+4.244693e+00*S37+5.513813e+01*S38+2.581070e+00*S39'
.param V17='V17_part4+3.157156e+00*S40+2.466713e+02*S41+1.857474e+00*S42+4.033303e+00*S43+2.219027e-02*S44'
.param V18_part1='(-8.429408e-01)*S0+(-1.973536e+00)*S1+(-1.327220e+00)*S2+(-1.714636e+00)*S3+(-1.485238e+00)*S4+(-2.807915e+00)*S5+(-5.498152e-01)*S6+(-1.390695e+00)*S7+(-1.324017e+00)*S8+(-1.314528e+00)*S9'
.param V18_part2='V18_part1+(-2.033006e+00)*S10+1.375497e+00*S11+(-7.066713e-01)*S12+(-1.872604e+00)*S13+(-2.021186e+00)*S14+(-1.027262e+00)*S15+(-2.594538e+00)*S16+(-1.447906e+00)*S17+(-3.009592e+00)*S18+(-2.467128e+00)*S19'
.param V18_part3='V18_part2+(-4.804727e+00)*S20+(-7.813596e-01)*S21+(-2.448961e+00)*S22+(-2.801138e+00)*S23+(-1.017703e+00)*S24+(-1.360841e+00)*S25+(-2.947402e+00)*S26+(-1.658121e+00)*S27+(-3.010829e+00)*S28+(-3.845838e+00)*S29'
.param V18_part4='V18_part3+(-1.400168e+00)*S30+(-2.480051e+00)*S31+(-3.303844e+00)*S32+(-4.371288e-01)*S33+(-3.385653e+00)*S34+(-5.513220e+00)*S35+(-2.035822e+00)*S36+0.000000e+00*S37+(-3.816660e+00)*S38+(-2.607351e+00)*S39'
.param V18='V18_part4+(-3.758561e+00)*S40+(-6.406162e+00)*S41+(-2.051831e+00)*S42+(-3.818135e+00)*S43+(-4.441254e+00)*S44'
.param V19_part1='6.147821e+00*S0+9.335217e+00*S1+5.482948e+00*S2+3.863602e+00*S3+3.260396e+00*S4+4.059460e+00*S5+6.401810e+00*S6+6.524141e+00*S7+7.061123e+00*S8+5.488003e+00*S9'
.param V19_part2='V19_part1+4.961205e+00*S10+1.733089e-01*S11+5.142948e+00*S12+5.653583e+00*S13+3.120531e+00*S14+7.803401e+00*S15+8.672487e+00*S16+5.370456e+00*S17+7.552421e+00*S18+5.795474e+00*S19'
.param V19_part3='V19_part2+7.997283e+00*S20+7.361309e+00*S21+7.459241e+00*S22+3.474705e+00*S23+5.766554e+00*S24+8.218757e-01*S25+6.498040e+00*S26+6.526617e+00*S27+7.475438e+00*S28+3.732586e+00*S29'
.param V19_part4='V19_part3+5.955123e+00*S30+7.002413e+00*S31+6.789640e+00*S32+4.320304e+00*S33+8.073309e+00*S34+9.845410e+00*S35+7.461035e+00*S36+0.000000e+00*S37+4.746199e+00*S38+8.059694e+00*S39'
.param V19='V19_part4+6.269870e+00*S40+1.084136e+01*S41+7.515931e+00*S42+8.952651e+00*S43+5.624833e+00*S44'
.param V20_part1='3.434186e+00*S0+3.974430e+00*S1+5.846811e+00*S2+6.361683e+00*S3+5.030221e+00*S4+6.775072e+00*S5+1.685299e+00*S6+3.057414e+00*S7+3.239446e+00*S8+2.605819e+00*S9'
.param V20_part2='V20_part1+3.750684e+00*S10+4.036001e+00*S11+6.215350e+00*S12+8.922429e+00*S13+8.028138e+00*S14+3.908098e+00*S15+5.246982e+00*S16+6.877648e+00*S17+7.381886e+00*S18+9.072982e+00*S19'
.param V20_part3='V20_part2+9.645918e+00*S20+6.636852e+00*S21+1.107989e+01*S22+1.219896e+01*S23+8.075152e+00*S24+7.666840e+00*S25+1.215826e+01*S26+1.188941e+01*S27+1.545833e+01*S28+1.362881e+01*S29'
.param V20_part4='V20_part3+1.054980e+01*S30+1.372041e+01*S31+1.676254e+01*S32+3.681273e+00*S33+1.891029e+01*S34+2.110513e+01*S35+1.295972e+01*S36+0.000000e+00*S37+1.115344e+01*S38+1.818935e+01*S39'
.param V20='V20_part4+1.316618e+01*S40+2.715615e+01*S41+1.555364e+01*S42+2.033942e+01*S43+1.219168e+01*S44'
.param V21_part1='7.641326e+00*S0+1.000000e+04*S1+7.003998e+00*S2+(-1.984136e+01)*S3+2.572968e-02*S4+(-1.555039e+01)*S5+4.475841e+01*S6+2.698357e+02*S7+7.934484e+03*S8+8.042099e+00*S9'
.param V21_part2='V21_part1+(-7.276629e+00)*S10+1.346275e+02*S11+8.311077e+00*S12+5.617932e+00*S13+4.326011e+03*S14+7.285048e+01*S15+7.049702e+01*S16+5.415058e+00*S17+4.984605e+00*S18+4.592060e+00*S19'
.param V21_part3='V21_part2+3.525154e+00*S20+1.633481e+02*S21+5.058414e+00*S22+2.957863e+00*S23+1.000000e+04*S24+2.899561e+01*S25+(-5.932573e+01)*S26+(-1.572099e+02)*S27+2.853790e+00*S28+2.356164e+00*S29'
.param V21_part4='V21_part3+3.688994e+00*S30+5.755149e+00*S31+3.927547e+00*S32+1.000000e+04*S33+9.455920e+00*S34+3.027768e+00*S35+(-1.511170e+03)*S36+(-1.213865e+01)*S37+1.181559e+03*S38+(-9.001255e+02)*S39'
.param V21='V21_part4+3.074290e+01*S40+3.592460e+00*S41+(-1.884089e+02)*S42+2.520508e+00*S43+7.008167e+00*S44'
.param V22_part1='(-2.530062e+00)*S0+(-4.182849e+01)*S1+(-5.470653e+00)*S2+(-8.949616e+00)*S3+(-2.569953e-01)*S4+4.290965e+00*S5+3.630977e+01*S6+(-3.252556e+00)*S7+4.905830e+02*S8+(-3.050141e+00)*S9'
.param V22_part2='V22_part1+6.864084e+00*S10+(-1.727736e+01)*S11+(-1.459312e+01)*S12+(-4.747788e+00)*S13+3.668134e+03*S14+(-2.958056e+01)*S15+(-1.176858e+02)*S16+(-4.663106e+00)*S17+(-3.475879e+00)*S18+(-2.257728e+00)*S19'
.param V22_part3='V22_part2+(-1.758787e+00)*S20+(-1.445747e+02)*S21+(-3.399611e+00)*S22+(-1.279075e+00)*S23+(-1.000000e+04)*S24+(-8.797900e+00)*S25+5.602647e+00*S26+1.104336e+03*S27+(-2.729335e+00)*S28+(-1.777435e+00)*S29'
.param V22_part4='V22_part3+(-6.380426e+00)*S30+(-4.416273e+00)*S31+(-2.330022e+00)*S32+(-9.330489e+00)*S33+(-8.650532e+00)*S34+(-1.950181e+00)*S35+1.000000e+04*S36+(-1.047554e+01)*S37+(-1.059983e+01)*S38+2.390742e+03*S39'
.param V22='V22_part4+(-1.131683e+02)*S40+(-1.987294e+00)*S41+(-1.548915e+03)*S42+(-1.638123e+00)*S43+(-2.979340e+00)*S44'
.param V23_part1='(-5.329096e+00)*S0+1.118624e+01*S1+(-1.116608e+00)*S2+8.187759e+01*S3+7.467650e+00*S4+3.817659e+01*S5+2.822876e+03*S6+(-2.156621e+02)*S7+(-8.585129e+03)*S8+(-2.549124e+00)*S9'
.param V23_part2='V23_part1+2.077969e+01*S10+(-1.051783e+02)*S11+3.212858e+00*S12+(-2.699510e-01)*S13+8.889644e+03*S14+(-4.119584e+01)*S15+7.663556e+00*S16+(-6.978763e-05)*S17+(-7.464549e-01)*S18+(-1.189910e+00)*S19'
.param V23_part3='V23_part2+(-2.646188e-01)*S20+(-9.693039e+01)*S21+(-9.223125e-01)*S22+(-6.483189e-01)*S23+1.000000e+04*S24+(-2.917937e+01)*S25+3.141581e+02*S26+6.182164e+01*S27+1.830224e+00*S28+4.797382e-01*S29'
.param V23_part4='V23_part3+1.776567e+00*S30+(-8.227082e-01)*S31+(-8.671410e-02)*S32+2.850780e-01*S33+1.058309e-01*S34+6.214853e-02*S35+4.987609e+02*S36+1.138311e+02*S37+(-2.189480e+03)*S38+2.860636e+03*S39'
.param V23='V23_part4+2.974445e+02*S40+(-3.006631e-01)*S41+4.431294e+03*S42+(-8.803214e-01)*S43+(-5.702795e+00)*S44'
.param V24_part1='1.289495e+01*S0+8.214366e+00*S1+5.935569e+00*S2+(-3.330953e+01)*S3+0.000000e+00*S4+(-3.269216e+00)*S5+1.730318e+01*S6+9.785570e+00*S7+0.000000e+00*S8+2.393123e+01*S9'
.param V24_part2='V24_part1+0.000000e+00*S10+4.568916e+01*S11+2.209369e+00*S12+0.000000e+00*S13+9.445085e+00*S14+5.368662e+00*S15+(-7.836725e-02)*S16+1.156848e+01*S17+1.476207e+01*S18+0.000000e+00*S19'
.param V24_part3='V24_part2+3.024305e+01*S20+8.319299e+00*S21+1.181197e+01*S22+0.000000e+00*S23+7.803198e+00*S24+(-1.588827e+01)*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V24_part4='V24_part3+0.000000e+00*S30+1.634205e+00*S31+7.431590e+01*S32+4.352058e+01*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+(-7.942523e+01)*S37+(-3.799134e+00)*S38+0.000000e+00*S39'
.param V24='V24_part4+(-7.368306e+01)*S40+8.641395e+01*S41+2.273829e+01*S42+0.000000e+00*S43+(-1.785952e+02)*S44'
.param V25_part1='2.573194e+01*S0+4.765803e+01*S1+7.243961e+01*S2+7.366235e+01*S3+0.000000e+00*S4+6.139426e+00*S5+2.881538e+01*S6+5.482533e+01*S7+0.000000e+00*S8+1.659104e+01*S9'
.param V25_part2='V25_part1+0.000000e+00*S10+(-6.663844e+01)*S11+9.672551e+01*S12+0.000000e+00*S13+(-7.920614e+00)*S14+4.845207e+01*S15+4.759683e+01*S16+6.180701e+01*S17+5.047493e+01*S18+0.000000e+00*S19'
.param V25_part3='V25_part2+3.424365e+01*S20+(-2.328612e+01)*S21+5.585503e+01*S22+0.000000e+00*S23+1.608383e+02*S24+1.778689e+01*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V25_part4='V25_part3+0.000000e+00*S30+6.485973e+01*S31+(-5.669820e+01)*S32+1.406869e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+3.086380e+02*S37+3.801481e+01*S38+0.000000e+00*S39'
.param V25='V25_part4+5.064014e+02*S40+(-8.884978e+00)*S41+(-2.403992e+01)*S42+0.000000e+00*S43+3.699237e+01*S44'
.param V26_part1='2.060222e+01*S0+1.512087e+01*S1+4.819005e+00*S2+1.438907e+01*S3+0.000000e+00*S4+4.266345e+01*S5+3.341929e+00*S6+1.766079e+01*S7+0.000000e+00*S8+(-7.344980e+00)*S9'
.param V26_part2='V26_part1+0.000000e+00*S10+4.754474e+01*S11+7.234712e+00*S12+0.000000e+00*S13+4.235236e+00*S14+2.430527e+01*S15+1.673450e+01*S16+1.047511e+01*S17+1.432559e+01*S18+0.000000e+00*S19'
.param V26_part3='V26_part2+1.282914e+01*S20+1.004864e+01*S21+2.616318e+01*S22+0.000000e+00*S23+3.576993e+01*S24+6.883704e+01*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V26_part4='V26_part3+0.000000e+00*S30+6.282989e+01*S31+1.177782e+02*S32+1.849870e+01*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+2.575791e+02*S37+4.270742e+02*S38+0.000000e+00*S39'
.param V26='V26_part4+3.548936e+02*S40+7.283208e+00*S41+1.857250e+02*S42+0.000000e+00*S43+1.220778e+03*S44'
.param V27_part1='(-7.446552e-01)*S0+(-1.898495e+00)*S1+(-1.407235e+00)*S2+(-1.541858e+00)*S3+(-1.317138e+00)*S4+(-2.661111e+00)*S5+(-5.571332e-01)*S6+(-1.370162e+00)*S7+(-1.317124e+00)*S8+(-1.279505e+00)*S9'
.param V27_part2='V27_part1+(-1.977743e+00)*S10+1.831187e+00*S11+(-7.305009e-01)*S12+(-1.930505e+00)*S13+(-1.965030e+00)*S14+(-1.030879e+00)*S15+(-2.570357e+00)*S16+(-1.447664e+00)*S17+(-3.003010e+00)*S18+(-2.284335e+00)*S19'
.param V27_part3='V27_part2+(-4.817454e+00)*S20+(-7.759026e-01)*S21+(-2.455169e+00)*S22+(-2.812212e+00)*S23+(-1.006930e+00)*S24+(-1.272493e+00)*S25+(-2.863084e+00)*S26+(-1.655032e+00)*S27+(-3.009326e+00)*S28+(-3.855967e+00)*S29'
.param V27_part4='V27_part3+(-1.405063e+00)*S30+(-2.557308e+00)*S31+(-3.711627e+00)*S32+(-4.370284e-01)*S33+(-3.048084e+00)*S34+(-5.514737e+00)*S35+(-2.031911e+00)*S36+0.000000e+00*S37+(-3.822303e+00)*S38+(-2.615100e+00)*S39'
.param V27='V27_part4+(-3.772131e+00)*S40+(-6.092393e+00)*S41+(-2.056510e+00)*S42+(-3.825760e+00)*S43+(-4.453765e+00)*S44'
.param V28_part1='5.079409e+00*S0+8.994092e+00*S1+5.930378e+00*S2+3.232759e+00*S3+3.033514e+00*S4+3.976925e+00*S5+6.389075e+00*S6+6.558447e+00*S7+7.056286e+00*S8+5.499262e+00*S9'
.param V28_part2='V28_part1+4.992806e+00*S10+(-4.933769e-01)*S11+5.577447e+00*S12+5.687176e+00*S13+3.018546e+00*S14+7.753917e+00*S15+8.654672e+00*S16+5.364085e+00*S17+7.602462e+00*S18+5.613408e+00*S19'
.param V28_part3='V28_part2+8.032672e+00*S20+7.273359e+00*S21+7.469938e+00*S22+3.480501e+00*S23+5.763883e+00*S24+9.039376e-01*S25+6.446420e+00*S26+6.530322e+00*S27+7.453737e+00*S28+3.739922e+00*S29'
.param V28_part4='V28_part3+5.969857e+00*S30+6.663421e+00*S31+7.187925e+00*S32+4.337568e+00*S33+7.866658e+00*S34+9.840766e+00*S35+7.470045e+00*S36+0.000000e+00*S37+4.749255e+00*S38+8.022768e+00*S39'
.param V28='V28_part4+6.295735e+00*S40+1.034639e+01*S41+7.553700e+00*S42+8.960689e+00*S43+5.638673e+00*S44'
.param V29_part1='3.650486e+00*S0+3.902679e+00*S1+5.789114e+00*S2+6.424189e+00*S3+5.269303e+00*S4+6.515474e+00*S5+1.590605e+00*S6+2.881591e+00*S7+3.072263e+00*S8+2.406439e+00*S9'
.param V29_part2='V29_part1+3.334839e+00*S10+3.941932e+00*S11+5.913793e+00*S12+8.912707e+00*S13+7.831093e+00*S14+3.836532e+00*S15+5.115418e+00*S16+6.823554e+00*S17+7.206177e+00*S18+8.869310e+00*S19'
.param V29_part3='V29_part2+9.499260e+00*S20+6.541347e+00*S21+1.093888e+01*S22+1.207117e+01*S23+7.776976e+00*S24+6.865066e+00*S25+1.189074e+01*S26+1.169818e+01*S27+1.534301e+01*S28+1.345980e+01*S29'
.param V29_part4='V29_part3+1.041781e+01*S30+1.386554e+01*S31+1.689209e+01*S32+3.488720e+00*S33+1.824339e+01*S34+2.096830e+01*S35+1.277348e+01*S36+0.000000e+00*S37+1.098021e+01*S38+1.804362e+01*S39'
.param V29='V29_part4+1.294998e+01*S40+2.742984e+01*S41+1.535597e+01*S42+2.019543e+01*S43+1.203031e+01*S44'
.param V30_part1='6.439307e+00*S0+8.595833e+00*S1+8.638807e+00*S2+4.515546e+00*S3+1.423750e+01*S4+5.905511e+00*S5+1.585245e+02*S6+5.626454e+00*S7+8.612888e+00*S8+8.451040e+00*S9'
.param V30_part2='V30_part1+6.225225e+00*S10+2.625133e+00*S11+1.469176e+01*S12+7.453185e+00*S13+1.583309e+01*S14+9.493998e+00*S15+5.157877e+01*S16+6.334700e+00*S17+4.950543e+00*S18+4.752686e+00*S19'
.param V30_part3='V30_part2+3.303442e+00*S20+1.028537e+01*S21+8.353408e+00*S22+2.282890e+03*S23+5.541823e+00*S24+(-4.263972e+01)*S25+3.509873e+00*S26+3.317537e+00*S27+8.539603e+00*S28+2.534996e+02*S29'
.param V30_part4='V30_part3+5.615675e+03*S30+5.761129e+00*S31+4.470812e+00*S32+4.263276e+00*S33+6.283993e+00*S34+2.596432e+00*S35+2.898480e+00*S36+3.862808e+00*S37+2.154144e+00*S38+3.137773e+03*S39'
.param V30='V30_part4+9.908141e+00*S40+3.919759e+00*S41+3.016761e+00*S42+(-1.990870e+03)*S43+2.692522e+00*S44'
.param V31_part1='(-5.296120e+00)*S0+(-1.634737e+00)*S1+(-5.093999e+00)*S2+(-3.489872e+00)*S3+(-1.056178e+01)*S4+(-2.482478e+00)*S5+2.545056e-03*S6+(-3.452594e+00)*S7+(-2.048613e+00)*S8+(-3.235871e+00)*S9'
.param V31_part2='V31_part1+(-3.127993e+00)*S10+(-4.997481e-01)*S11+(-1.549662e+01)*S12+(-5.385927e+00)*S13+(-7.759956e+00)*S14+(-3.838980e+00)*S15+(-8.255268e+01)*S16+(-5.646917e+00)*S17+(-4.174527e+00)*S18+(-2.547878e+00)*S19'
.param V31_part3='V31_part2+(-1.899882e+00)*S20+(-9.301736e+00)*S21+(-5.339616e+00)*S22+1.000000e+04*S23+(-7.575829e+00)*S24+(-1.513711e+01)*S25+(-1.820719e+00)*S26+(-5.327330e+00)*S27+(-8.570120e+00)*S28+(-7.384239e+00)*S29'
.param V31_part4='V31_part3+(-1.200624e+02)*S30+(-4.672625e+00)*S31+(-2.487445e+00)*S32+(-4.570073e+00)*S33+(-3.337197e+00)*S34+2.141973e+00*S35+(-4.511997e+00)*S36+(-3.448181e+00)*S37+(-1.767162e+00)*S38+1.119225e+00*S39'
.param V31='V31_part4+(-5.566055e+00)*S40+(-8.036476e+00)*S41+(-4.279537e+00)*S42+(-2.074636e+00)*S43+(-2.537981e+00)*S44'
.param V32_part1='(-1.606316e+00)*S0+(-4.447808e+00)*S1+(-3.299570e+00)*S2+5.256348e-01*S3+(-8.929378e-01)*S4+(-9.562814e-01)*S5+(-1.375075e+02)*S6+(-1.865218e+00)*S7+(-6.701102e+00)*S8+(-2.615187e+00)*S9'
.param V32_part2='V32_part1+(-1.835387e+00)*S10+8.926968e-01*S11+(-9.006592e+00)*S12+(-2.696540e+00)*S13+(-3.807237e+00)*S14+(-6.939285e+00)*S15+4.723096e+00*S16+(-1.232185e-01)*S17+5.738261e-01*S18+(-1.011798e+00)*S19'
.param V32_part3='V32_part2+2.985940e-01*S20+(-6.879052e+00)*S21+(-3.531070e+00)*S22+(-4.070641e+03)*S23+(-1.141538e+00)*S24+3.197105e+02*S25+(-3.527516e-02)*S26+1.286089e+00*S27+1.261938e+00*S28+(-4.507402e+02)*S29'
.param V32_part4='V32_part3+4.643228e+01*S30+(-7.645335e-01)*S31+(-6.706995e-01)*S32+(-1.986222e+00)*S33+(-4.552872e+00)*S34+(-3.603694e+00)*S35+1.132179e+00*S36+(-3.890717e-01)*S37+7.117685e-01*S38+(-5.866465e+03)*S39'
.param V32='V32_part4+(-8.867978e+00)*S40+3.599480e+01*S41+3.634733e-01*S42+9.992032e+03*S43+2.302293e+00*S44'
.param V33_part1='2.740831e+01*S0+6.357699e+00*S1+3.560445e+00*S2+2.235792e+01*S3+(-1.572010e+01)*S4+1.162716e+01*S5+0.000000e+00*S6+8.362758e+00*S7+(-8.617378e-01)*S8+2.382696e+01*S9'
.param V33_part2='V33_part1+3.337918e+00*S10+6.641633e+01*S11+4.676240e+00*S12+(-4.142600e+01)*S13+0.000000e+00*S14+4.796291e+00*S15+(-7.680713e-01)*S16+0.000000e+00*S17+0.000000e+00*S18+2.064109e+01*S19'
.param V33_part3='V33_part2+1.925905e+01*S20+6.075910e+00*S21+1.257366e+01*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+6.163247e+01*S26+0.000000e+00*S27+(-2.136656e+00)*S28+0.000000e+00*S29'
.param V33_part4='V33_part3+0.000000e+00*S30+2.075338e+01*S31+3.358914e+01*S32+(-4.512449e+01)*S33+5.266034e+01*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V33='V33_part4+0.000000e+00*S40+5.729913e+00*S41+0.000000e+00*S42+(-7.233191e-01)*S43+0.000000e+00*S44'
.param V34_part1='1.569445e+01*S0+5.078397e+01*S1+6.105005e+01*S2+1.687882e+01*S3+1.444517e+02*S4+2.778777e+01*S5+0.000000e+00*S6+5.423467e+01*S7+5.165081e+01*S8+1.495400e+01*S9'
.param V34_part2='V34_part1+5.829504e+01*S10+(-2.702217e+01)*S11+5.435651e+01*S12+9.857913e+01*S13+0.000000e+00*S14+4.934860e+01*S15+4.759431e+01*S16+0.000000e+00*S17+0.000000e+00*S18+5.344506e+01*S19'
.param V34_part3='V34_part2+4.650969e+01*S20+6.816473e+01*S21+5.552902e+01*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+(-9.013685e+00)*S26+0.000000e+00*S27+(-1.742796e+00)*S28+0.000000e+00*S29'
.param V34_part4='V34_part3+0.000000e+00*S30+7.188731e-01*S31+(-9.148462e+00)*S32+1.121298e+02*S33+(-1.513768e+02)*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V34='V34_part4+0.000000e+00*S40+(-9.987437e+01)*S41+0.000000e+00*S42+(-5.676854e+01)*S43+0.000000e+00*S44'
.param V35_part1='(-7.499671e-01)*S0+1.517837e+01*S1+1.291585e+01*S2+1.380924e+01*S3+4.902977e+01*S4+1.345710e+01*S5+0.000000e+00*S6+1.842696e+01*S7+3.189284e+01*S8+(-7.603797e+00)*S9'
.param V35_part2='V35_part1+(-2.531970e+00)*S10+(-5.527724e+00)*S11+2.221167e+01*S12+1.034603e+02*S13+0.000000e+00*S14+2.384149e+01*S15+1.681393e+01*S16+0.000000e+00*S17+0.000000e+00*S18+1.142946e+01*S19'
.param V35_part3='V35_part2+1.861880e+01*S20+2.136142e+01*S21+2.430987e+01*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+2.358436e+01*S26+0.000000e+00*S27+2.637349e+02*S28+0.000000e+00*S29'
.param V35_part4='V35_part3+0.000000e+00*S30+8.132437e+01*S31+1.301676e+02*S32+1.443021e+02*S33+3.323190e+02*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V35='V35_part4+0.000000e+00*S40+4.676762e+02*S41+0.000000e+00*S42+4.107849e+02*S43+0.000000e+00*S44'
.param V36_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-3.592197e+00)*S3+(-1.690971e+00)*S4+(-3.030483e+00)*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+(-1.666108e+00)*S9'
.param V36_part2='V36_part1+(-3.223262e-01)*S10+(-9.059403e+00)*S11+0.000000e+00*S12+0.000000e+00*S13+(-1.500423e+00)*S14+0.000000e+00*S15+1.704838e-01*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V36_part3='V36_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+(-1.613283e+00)*S23+0.000000e+00*S24+(-1.695539e+00)*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+3.484314e-01*S29'
.param V36_part4='V36_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+(-3.171850e+00)*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+(-5.024756e+00)*S37+(-2.971133e-01)*S38+0.000000e+00*S39'
.param V36='V36_part4+7.874245e-01*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+(-7.753793e-01)*S44'
.param V37_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+7.625995e+00*S3+3.760998e+00*S4+6.418083e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+3.370982e+00*S9'
.param V37_part2='V37_part1+9.968283e-01*S10+1.217653e+01*S11+0.000000e+00*S12+0.000000e+00*S13+5.745960e+00*S14+0.000000e+00*S15+8.176525e-01*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V37_part3='V37_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+1.058702e+01*S23+0.000000e+00*S24+1.104054e+01*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+6.090249e+00*S29'
.param V37_part4='V37_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+6.352589e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+1.299258e+01*S37+5.133098e+00*S38+0.000000e+00*S39'
.param V37='V37_part4+5.047695e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+5.489162e+00*S44'
.param V38_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+9.243619e-01*S3+6.295844e+00*S4+3.267139e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+2.426574e+00*S9'
.param V38_part2='V38_part1+3.558918e+00*S10+3.638779e+00*S11+0.000000e+00*S12+0.000000e+00*S13+5.894534e+00*S14+0.000000e+00*S15+5.074234e-01*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V38_part3='V38_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+8.577806e-01*S23+0.000000e+00*S24+5.344147e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+1.190809e+01*S29'
.param V38_part4='V38_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+2.106570e+01*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+3.486739e+01*S37+1.900057e+01*S38+0.000000e+00*S39'
.param V38='V38_part4+1.667227e+01*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+2.503979e+01*S44'
.param V39_part1='0.000000e+00*S0+0.000000e+00*S1+1.000000e+04*S2+5.756377e+00*S3+9.933750e+00*S4+3.996054e+00*S5+0.000000e+00*S6+5.406923e+00*S7+8.744584e+00*S8+2.905985e+00*S9'
.param V39_part2='V39_part1+5.582513e+00*S10+2.414146e+00*S11+1.272855e+03*S12+(-1.956746e+02)*S13+0.000000e+00*S14+0.000000e+00*S15+1.370826e+00*S16+(-3.583406e+01)*S17+6.161758e+01*S18+(-3.010533e+02)*S19'
.param V39_part3='V39_part2+1.676813e+02*S20+1.035715e+01*S21+1.048997e+01*S22+7.241776e+02*S23+1.000000e+04*S24+4.009159e+00*S25+4.488869e+00*S26+1.175993e+03*S27+4.815910e+03*S28+(-9.851905e+01)*S29'
.param V39_part4='V39_part3+2.314144e+02*S30+(-3.169260e+02)*S31+(-3.093418e+01)*S32+(-1.989916e+03)*S33+5.094621e+00*S34+4.454373e+01*S35+5.345776e+03*S36+8.125002e+01*S37+1.000000e+04*S38+2.804420e+00*S39'
.param V39='V39_part4+5.781016e+00*S40+0.000000e+00*S41+2.602668e+02*S42+(-5.133616e+01)*S43+1.923381e+03*S44'
.param V40_part1='0.000000e+00*S0+0.000000e+00*S1+(-4.054794e+03)*S2+(-3.858478e+00)*S3+(-5.140427e+00)*S4+(-2.103741e+00)*S5+0.000000e+00*S6+(-3.584918e+00)*S7+(-2.390644e+00)*S8+(-3.616249e+00)*S9'
.param V40_part2='V40_part1+(-2.613695e+00)*S10+(-7.834297e-01)*S11+(-7.421684e+00)*S12+(-2.054168e+00)*S13+0.000000e+00*S14+0.000000e+00*S15+(-3.405830e+00)*S16+(-7.336018e+01)*S17+(-1.569347e+01)*S18+7.771900e+00*S19'
.param V40_part3='V40_part2+(-4.869894e+00)*S20+(-7.561041e+00)*S21+(-9.110029e+00)*S22+(-2.639814e+00)*S23+(-1.000000e+04)*S24+(-3.081730e+00)*S25+(-2.132792e+00)*S26+(-2.466337e+01)*S27+(-7.267865e+00)*S28+(-6.902510e+00)*S29'
.param V40_part4='V40_part3+(-3.231660e+01)*S30+1.984795e+01*S31+2.580338e+01*S32+(-1.168920e+01)*S33+(-6.871923e+00)*S34+(-2.611193e+01)*S35+(-1.411784e+01)*S36+(-2.016220e+01)*S37+9.568000e+03*S38+(-3.821610e+00)*S39'
.param V40='V40_part4+(-5.887650e+00)*S40+0.000000e+00*S41+(-1.565000e-01)*S42+(-1.088166e+03)*S43+(-7.958755e-01)*S44'
.param V41_part1='0.000000e+00*S0+0.000000e+00*S1+(-4.957985e+03)*S2+(-1.143351e+00)*S3+(-4.742594e+00)*S4+(-5.523326e-01)*S5+0.000000e+00*S6+(-1.621453e+00)*S7+(-6.389988e+00)*S8+6.977452e-01*S9'
.param V41_part2='V41_part1+(-2.507007e+00)*S10+(-5.262803e-01)*S11+(-2.348131e+03)*S12+1.002162e+03*S13+0.000000e+00*S14+0.000000e+00*S15+1.392521e-01*S16+5.212190e+02*S17+(-4.466171e+01)*S18+1.493338e+03*S19'
.param V41_part3='V41_part2+(-1.533426e+02)*S20+(-8.252245e+00)*S21+1.167311e+01*S22+(-1.344981e+03)*S23+1.000000e+04*S24+(-6.103737e-01)*S25+(-1.680454e+00)*S26+(-2.173734e+03)*S27+(-9.007739e+03)*S28+5.615520e+02*S29'
.param V41_part4='V41_part3+(-3.987253e+02)*S30+1.586415e+03*S31+1.002827e+02*S32+1.000000e+04*S33+1.196678e+01*S34+(-9.113196e+00)*S35+(-1.000000e+04)*S36+(-1.134416e+02)*S37+5.971044e+03*S38+2.314158e-01*S39'
.param V41='V41_part4+(-9.411530e-01)*S40+0.000000e+00*S41+(-4.743013e+02)*S42+4.733998e+03*S43+3.607705e+00*S44'
.param V42_part1='4.802157e+03*S0+0.000000e+00*S1+0.000000e+00*S2+3.262500e+01*S3+0.000000e+00*S4+1.065662e+01*S5+0.000000e+00*S6+0.000000e+00*S7+2.337014e+00*S8+(-1.097177e+02)*S9'
.param V42_part2='V42_part1+2.325303e+01*S10+(-6.802326e+01)*S11+0.000000e+00*S12+5.775839e+01*S13+3.727426e+03*S14+7.667964e+02*S15+1.153920e+01*S16+9.911108e+00*S17+1.151736e+01*S18+1.656995e+01*S19'
.param V42_part3='V42_part2+0.000000e+00*S20+(-2.762497e+00)*S21+0.000000e+00*S22+(-1.224066e+01)*S23+0.000000e+00*S24+4.746542e+00*S25+5.295753e+01*S26+1.935671e+01*S27+0.000000e+00*S28+3.777038e+01*S29'
.param V42_part4='V42_part3+1.456626e+01*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+7.617514e+00*S36+0.000000e+00*S37+(-1.397037e+02)*S38+2.837966e+00*S39'
.param V42='V42_part4+(-2.634450e+01)*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V43_part1='4.802157e+03*S0+0.000000e+00*S1+0.000000e+00*S2+1.603739e+01*S3+0.000000e+00*S4+8.121287e+01*S5+0.000000e+00*S6+0.000000e+00*S7+5.688505e+01*S8+1.643551e+02*S9'
.param V43_part2='V43_part1+7.526312e+01*S10+2.131059e+02*S11+0.000000e+00*S12+(-1.403076e+01)*S13+3.215509e+03*S14+(-5.418263e+01)*S15+3.215957e+02*S16+6.842298e+01*S17+5.862496e+01*S18+5.573919e+01*S19'
.param V43_part3='V43_part2+0.000000e+00*S20+9.601390e+01*S21+0.000000e+00*S22+3.688326e+01*S23+0.000000e+00*S24+2.135339e+02*S25+1.161660e+00*S26+6.315262e+01*S27+0.000000e+00*S28+2.876419e+01*S29'
.param V43_part4='V43_part3+1.234148e+02*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+5.711395e+01*S36+0.000000e+00*S37+1.495759e+02*S38+(-1.115094e+02)*S39'
.param V43='V43_part4+6.143888e+01*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V44_part1='4.802157e+03*S0+0.000000e+00*S1+0.000000e+00*S2+(-4.633892e+00)*S3+0.000000e+00*S4+(-3.273545e+01)*S5+0.000000e+00*S6+0.000000e+00*S7+2.411623e+01*S8+1.285639e+02*S9'
.param V44_part2='V44_part1+1.736226e+00*S10+(-3.678926e+01)*S11+0.000000e+00*S12+(-3.256880e+01)*S13+3.464113e+03*S14+2.870539e+02*S15+2.036703e+01*S16+6.802599e+00*S17+1.605945e+01*S18+1.671523e+01*S19'
.param V44_part3='V44_part2+0.000000e+00*S20+1.451844e+01*S21+0.000000e+00*S22+3.749975e+02*S23+0.000000e+00*S24+(-5.282725e+01)*S25+3.111969e+01*S26+9.999333e+01*S27+0.000000e+00*S28+4.139851e+02*S29'
.param V44_part4='V44_part3+7.106405e+01*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+1.473988e+02*S36+0.000000e+00*S37+2.894530e+02*S38+2.905352e+02*S39'
.param V44='V44_part4+2.465327e+01*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V45_part1='(-1.415109e+00)*S0+9.417308e+03*S1+1.000000e+04*S2+5.640645e+00*S3+9.998305e-01*S4+6.871015e+00*S5+5.200642e-01*S6+8.265502e+02*S7+6.940305e+00*S8+1.657305e+02*S9'
.param V45_part2='V45_part1+9.278796e+03*S10+3.136395e+01*S11+(-7.922633e+00)*S12+3.965768e-01*S13+(-1.111873e+01)*S14+2.052816e+01*S15+1.000000e+04*S16+1.281660e+01*S17+6.356241e+00*S18+9.569634e+01*S19'
.param V45_part3='V45_part2+7.672674e+01*S20+3.779692e+01*S21+6.931796e+01*S22+0.000000e+00*S23+1.726228e+02*S24+(-2.617233e+01)*S25+1.575192e+01*S26+0.000000e+00*S27+1.000000e+04*S28+0.000000e+00*S29'
.param V45_part4='V45_part3+0.000000e+00*S30+1.000000e+04*S31+5.131763e+02*S32+6.912246e+01*S33+(-4.088622e+01)*S34+5.612507e+01*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V45='V45_part4+8.117503e+00*S40+1.218554e+01*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V46_part1='1.257130e+02*S0+5.698090e+02*S1+1.000000e+04*S2+(-9.686072e-01)*S3+(-8.028480e-01)*S4+(-9.257856e-02)*S5+(-1.279635e+00)*S6+7.908653e+01*S7+(-3.283346e+00)*S8+1.215638e+02*S9'
.param V46_part2='V46_part1+1.000000e+04*S10+5.797996e+00*S11+8.217634e+01*S12+(-5.168563e-01)*S13+9.128729e+01*S14+(-5.398925e+01)*S15+1.000000e+04*S16+2.756359e+00*S17+7.877166e-01*S18+1.936003e+02*S19'
.param V46_part3='V46_part2+(-1.356836e+02)*S20+(-1.708387e+02)*S21+(-1.735561e+03)*S22+0.000000e+00*S23+8.421886e+02*S24+1.256933e+03*S25+(-3.151842e-01)*S26+0.000000e+00*S27+1.000000e+04*S28+0.000000e+00*S29'
.param V46_part4='V46_part3+0.000000e+00*S30+1.000000e+04*S31+1.000000e+04*S32+4.754230e+00*S33+2.844005e+01*S34+8.520415e+03*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V46='V46_part4+2.105373e+01*S40+1.269796e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V47_part1='(-3.251459e+01)*S0+7.994881e+02*S1+(-6.166480e+03)*S2+(-3.461221e+00)*S3+1.036636e-01*S4+(-5.676036e+00)*S5+1.376200e-01*S6+2.990368e+03*S7+(-3.068983e+00)*S8+(-1.785825e+02)*S9'
.param V47_part2='V47_part1+(-1.715675e+01)*S10+(-2.821925e+01)*S11+(-1.756519e+01)*S12+2.144836e-01*S13+(-9.925024e+01)*S14+4.662721e+01*S15+1.000000e+04*S16+(-1.666471e+01)*S17+(-5.631802e+00)*S18+(-2.554977e+02)*S19'
.param V47_part3='V47_part2+9.908405e+01*S20+1.712464e+02*S21+5.803861e+03*S22+0.000000e+00*S23+6.607789e+02*S24+(-9.310664e+02)*S25+(-2.810186e+01)*S26+0.000000e+00*S27+1.000000e+04*S28+0.000000e+00*S29'
.param V47_part4='V47_part3+0.000000e+00*S30+1.000000e+04*S31+6.151144e+01*S32+6.329869e+01*S33+1.697259e+02*S34+6.668003e+03*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V47='V47_part4+1.556641e+01*S40+(-2.352929e+01)*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V48_part1='(-1.552368e-01)*S0+(-2.649492e-01)*S1+(-4.735998e-01)*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+(-2.270623e-01)*S9'
.param V48_part2='V48_part1+0.000000e+00*S10+3.909301e-01*S11+(-3.630081e-01)*S12+0.000000e+00*S13+1.252796e+00*S14+(-2.106542e-01)*S15+(-1.977283e-01)*S16+(-7.312463e-01)*S17+0.000000e+00*S18+(-1.498590e+00)*S19'
.param V48_part3='V48_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+(-7.576875e-01)*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V48_part4='V48_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+(-2.916172e+01)*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V48='V48_part4+9.063599e+01*S40+(-4.342142e+01)*S41+0.000000e+00*S42+1.000000e+04*S43+0.000000e+00*S44'
.param V49_part1='5.711659e-01*S0+1.046422e+00*S1+1.304414e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+5.101255e-01*S9'
.param V49_part2='V49_part1+0.000000e+00*S10+(-1.413012e-01)*S11+3.294518e+00*S12+0.000000e+00*S13+(-5.960633e-01)*S14+1.102459e+00*S15+6.635872e-01*S16+3.025950e+00*S17+0.000000e+00*S18+2.052548e+00*S19'
.param V49_part3='V49_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+1.337021e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V49_part4='V49_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+5.278482e+01*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V49='V49_part4+4.448495e+00*S40+9.639351e+01*S41+0.000000e+00*S42+1.000000e+04*S43+0.000000e+00*S44'
.param V50_part1='3.530513e-01*S0+1.625078e-01*S1+2.328742e-01*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+1.752448e-01*S9'
.param V50_part2='V50_part1+0.000000e+00*S10+3.287675e-01*S11+8.758915e-01*S12+0.000000e+00*S13+(-7.162517e-02)*S14+1.878865e-01*S15+3.278864e-01*S16+7.594785e-01*S17+0.000000e+00*S18+1.352124e+00*S19'
.param V50_part3='V50_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+3.168359e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V50_part4='V50_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+3.501673e+01*S34+0.000000e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V50='V50_part4+(-7.105456e+00)*S40+(-4.444899e+01)*S41+0.000000e+00*S42+1.000000e+04*S43+0.000000e+00*S44'
.param V51_part1='1.446964e+00*S0+6.522860e+00*S1+0.000000e+00*S2+0.000000e+00*S3+8.727907e+00*S4+2.294294e+01*S5+5.207862e+00*S6+0.000000e+00*S7+0.000000e+00*S8+(-1.872729e+03)*S9'
.param V51_part2='V51_part1+3.058461e-02*S10+(-1.331352e-01)*S11+0.000000e+00*S12+0.000000e+00*S13+1.568942e+01*S14+9.910854e+00*S15+6.175925e+00*S16+3.159414e+00*S17+3.603206e+00*S18+0.000000e+00*S19'
.param V51_part3='V51_part2+4.290059e+00*S20+0.000000e+00*S21+5.787858e+00*S22+4.479741e+03*S23+0.000000e+00*S24+1.000000e+04*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V51_part4='V51_part3+1.098005e+03*S30+1.000000e+04*S31+1.000000e+04*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+1.000000e+04*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V51='V51_part4+0.000000e+00*S40+3.842008e+01*S41+4.617642e+03*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V52_part1='(-3.948858e+02)*S0+(-2.432204e+00)*S1+0.000000e+00*S2+0.000000e+00*S3+2.524242e+00*S4+2.748854e+01*S5+(-1.114502e+00)*S6+0.000000e+00*S7+0.000000e+00*S8+1.000000e+04*S9'
.param V52_part2='V52_part1+4.713955e-03*S10+(-6.971016e-02)*S11+0.000000e+00*S12+0.000000e+00*S13+(-5.835704e+00)*S14+(-2.891104e+00)*S15+3.044386e+00*S16+(-6.273656e+00)*S17+(-4.085200e+00)*S18+0.000000e+00*S19'
.param V52_part3='V52_part2+4.536418e-01*S20+0.000000e+00*S21+1.884610e+02*S22+4.785111e+03*S23+0.000000e+00*S24+1.000000e+04*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V52_part4='V52_part3+5.578035e+03*S30+1.000000e+04*S31+1.000000e+04*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+9.080540e+02*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V52='V52_part4+0.000000e+00*S40+(-1.473650e+01)*S41+7.103505e+02*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V53_part1='3.851302e+03*S0+(-2.722185e+00)*S1+0.000000e+00*S2+0.000000e+00*S3+(-1.030687e+01)*S4+1.147948e+01*S5+(-4.324999e+00)*S6+0.000000e+00*S7+0.000000e+00*S8+(-2.087937e+03)*S9'
.param V53_part2='V53_part1+(-7.303426e-04)*S10+1.032711e+00*S11+0.000000e+00*S12+0.000000e+00*S13+(-8.682046e+00)*S14+(-7.991307e+00)*S15+(-4.345982e+00)*S16+7.437906e+00*S17+3.943359e-01*S18+0.000000e+00*S19'
.param V53_part3='V53_part2+(-4.251185e+00)*S20+0.000000e+00*S21+(-1.407447e+02)*S22+1.000000e+04*S23+0.000000e+00*S24+1.727385e+03*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V53_part4='V53_part3+1.000000e+04*S30+1.000000e+04*S31+5.171578e+02*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+1.000000e+04*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V53='V53_part4+0.000000e+00*S40+4.338606e-01*S41+2.549420e+02*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V54_part1='0.000000e+00*S0+0.000000e+00*S1+1.000000e+04*S2+0.000000e+00*S3+0.000000e+00*S4+8.789371e+02*S5+0.000000e+00*S6+(-1.458981e+03)*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V54_part2='V54_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+(-1.875000e+00)*S18+0.000000e+00*S19'
.param V54_part3='V54_part2+(-5.929965e+00)*S20+6.626419e+00*S21+(-6.465168e-01)*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V54_part4='V54_part3+0.000000e+00*S30+(-5.238467e-01)*S31+(-1.237797e+00)*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+(-5.726726e+00)*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V54='V54_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V55_part1='0.000000e+00*S0+0.000000e+00*S1+1.000000e+04*S2+0.000000e+00*S3+0.000000e+00*S4+3.248454e+02*S5+0.000000e+00*S6+(-3.835033e+03)*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V55_part2='V55_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+5.116841e+00*S18+0.000000e+00*S19'
.param V55_part3='V55_part2+9.339735e+00*S20+5.705166e+01*S21+1.282366e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V55_part4='V55_part3+0.000000e+00*S30+1.829781e+00*S31+3.050123e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+2.684927e+01*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V55='V55_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V56_part1='0.000000e+00*S0+0.000000e+00*S1+1.000000e+04*S2+0.000000e+00*S3+0.000000e+00*S4+5.571058e+02*S5+0.000000e+00*S6+5.921843e+03*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V56_part2='V56_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+1.961465e+00*S18+0.000000e+00*S19'
.param V56_part3='V56_part2+3.850637e+00*S20+5.576023e-01*S21+1.563412e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V56_part4='V56_part3+0.000000e+00*S30+2.167580e-01*S31+1.146051e-01*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36+6.874775e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V56='V56_part4+0.000000e+00*S40+0.000000e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V57_part1='(-5.954281e+01)*S0+3.714225e+01*S1+5.527824e+01*S2+2.271384e+02*S3+0.000000e+00*S4+1.176746e+01*S5+2.429582e+01*S6+(-1.395390e+01)*S7+(-2.192693e+01)*S8+(-2.722101e+03)*S9'
.param V57_part2='V57_part1+(-1.999451e+03)*S10+(-2.904145e+01)*S11+8.761616e+01*S12+4.309317e+03*S13+6.166366e+02*S14+1.442579e+02*S15+6.863320e+00*S16+0.000000e+00*S17+0.000000e+00*S18+(-1.999049e+03)*S19'
.param V57_part3='V57_part2+2.545483e-01*S20+7.423597e+00*S21+0.000000e+00*S22+8.453754e+03*S23+0.000000e+00*S24+0.000000e+00*S25+9.401257e+03*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V57_part4='V57_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+3.262875e+00*S34+0.000000e+00*S35+0.000000e+00*S36+1.000000e+04*S37+0.000000e+00*S38+6.250000e+02*S39'
.param V57='V57_part4+9.201993e+01*S40+6.359028e+00*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V58_part1='2.149333e+01*S0+(-6.044472e+01)*S1+8.788213e+02*S2+1.299762e+01*S3+0.000000e+00*S4+(-1.901728e+01)*S5+(-2.124112e+00)*S6+2.574021e+02*S7+(-3.321460e-01)*S8+1.000000e+04*S9'
.param V58_part2='V58_part1+(-3.564103e-01)*S10+6.412175e+01*S11+(-9.841597e+00)*S12+(-6.431167e+02)*S13+6.459446e+00*S14+2.848688e+02*S15+3.338441e+00*S16+0.000000e+00*S17+0.000000e+00*S18+(-7.144356e-01)*S19'
.param V58_part3='V58_part2+2.305908e-01*S20+7.657927e+01*S21+0.000000e+00*S22+9.042868e+03*S23+0.000000e+00*S24+0.000000e+00*S25+(-1.000000e+04)*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V58_part4='V58_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+1.507075e+01*S34+0.000000e+00*S35+0.000000e+00*S36+1.000000e+04*S37+0.000000e+00*S38+1.000000e+04*S39'
.param V58='V58_part4+1.163439e+02*S40+(-1.389089e+00)*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V59_part1='3.226416e+02*S0+5.975747e+00*S1+(-3.664294e+02)*S2+1.126762e+02*S3+0.000000e+00*S4+1.353644e+01*S5+(-1.982038e+01)*S6+(-4.282699e+01)*S7+1.109238e+02*S8+3.556887e+01*S9'
.param V59_part2='V59_part1+1.000000e+04*S10+1.111488e+00*S11+(-1.515542e+02)*S12+(-6.942755e+03)*S13+(-1.081189e+03)*S14+(-2.381878e+02)*S15+(-4.926029e+00)*S16+0.000000e+00*S17+0.000000e+00*S18+1.000000e+04*S19'
.param V59_part3='V59_part2+(-4.051249e-01)*S20+(-4.309490e+01)*S21+0.000000e+00*S22+9.562975e+03*S23+0.000000e+00*S24+0.000000e+00*S25+2.997668e+03*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V59_part4='V59_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+(-1.821572e+01)*S34+0.000000e+00*S35+0.000000e+00*S36+1.000000e+04*S37+0.000000e+00*S38+1.000000e+04*S39'
.param V59='V59_part4+6.434488e+01*S40+(-6.159902e+00)*S41+0.000000e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V60_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-7.195321e-01)*S3+1.337438e+01*S4+(-1.405769e+00)*S5+3.745920e-02*S6+(-3.428705e-01)*S7+(-7.839102e-01)*S8+0.000000e+00*S9'
.param V60_part2='V60_part1+(-6.917994e-01)*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+2.698442e+02*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V60_part3='V60_part2+0.000000e+00*S20+(-5.174494e-01)*S21+0.000000e+00*S22+1.345850e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V60_part4='V60_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+7.648113e+03*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V60='V60_part4+1.037483e+02*S40+0.000000e+00*S41+5.723272e+02*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V61_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+1.664261e+00*S3+1.024852e+02*S4+1.810818e+00*S5+6.966115e-01*S6+1.026515e+00*S7+2.582100e+00*S8+0.000000e+00*S9'
.param V61_part2='V61_part1+9.215648e-01*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+6.131186e+02*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V61_part3='V61_part2+0.000000e+00*S20+1.478919e+00*S21+0.000000e+00*S22+(-1.717750e+00)*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V61_part4='V61_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+5.189756e+00*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V61='V61_part4+1.857614e+01*S40+0.000000e+00*S41+3.371642e+00*S42+0.000000e+00*S43+0.000000e+00*S44'
.param V62_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+1.268637e+00*S3+1.065370e+02*S4+1.626645e+00*S5+1.696771e-01*S6+2.038003e-01*S7+4.408709e-01*S8+0.000000e+00*S9'
.param V62_part2='V62_part1+4.064928e-01*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+1.000000e+04*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V62_part3='V62_part2+0.000000e+00*S20+1.645763e+00*S21+0.000000e+00*S22+4.680795e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V62_part4='V62_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+1.000000e+04*S35+0.000000e+00*S36+0.000000e+00*S37+0.000000e+00*S38+0.000000e+00*S39'
.param V62='V62_part4+(-9.788055e-01)*S40+0.000000e+00*S41+1.000000e+04*S42+0.000000e+00*S43+0.000000e+00*S44'
.param _P0='V0+V1*radius_+V2*w_'
.param _P1='0.5*(_P0+sqrt(_P0*_P0+0.001))'
.param _P2='1e-15*_P1'
.param _P3='V3+V4*radius_+V5/w_'
.param _P4='0.5*(_P3+sqrt(_P3*_P3+0.001))'
.param _P5='V6+V7*radius_+V8*w_'
.param _P6='0.5*(_P5+sqrt(_P5*_P5+0.001))'
.param _P7='1e-09*_P6'
.param _P8='1e-09*_P6'
.param _P9='V9+V10*radius_+V11/w_'
.param _P10='0.5*(_P9+sqrt(_P9*_P9+0.001))'
.param _P11='V12+V13*radius_+V14*w_'
.param _P12='0.5*(_P11+sqrt(_P11*_P11+0.001))'
.param _P13='1e-09*_P12'
.param _P14='V15+V16*radius_+V17*w_'
.param _P15='0.5*(atan(2*_P14)/1.5708+1)'
.param _P16='0.7064*_P15'
.param _P17='0.7064*_P15'
.param _P18='V18+V19*radius_+V20*w_'
.param _P19='0.5*(_P18+sqrt(_P18*_P18+0.001))'
.param _P20='V21+V22*radius_+V23*w_'
.param _P21='0.5*(_P20+sqrt(_P20*_P20+0.001))'
.param _P22='V24+V25*radius_+V26*w_'
.param _P23='0.5*(_P22+sqrt(_P22*_P22+0.001))'
.param _P24='V27+V28*radius_+V29*w_'
.param _P25='0.5*(_P24+sqrt(_P24*_P24+0.001))'
.param _P26='V30+V31*radius_+V32*w_'
.param _P27='0.5*(_P26+sqrt(_P26*_P26+0.001))'
.param _P28='V33+V34*radius_+V35*w_'
.param _P29='0.5*(_P28+sqrt(_P28*_P28+0.001))'
.param _P30='V36+V37*radius_+V38*w_'
.param _P31='0.5*(_P30+sqrt(_P30*_P30+0.001))'
.param _P32='V39+V40*radius_+V41*w_'
.param _P33='0.5*(_P32+sqrt(_P32*_P32+0.001))'
.param _P34='V42+V43*radius_+V44*w_'
.param _P35='0.5*(_P34+sqrt(_P34*_P34+0.001))'
.param _P36='1e-14*_P19'
.param _P37='100*_P21'
.param _P38='1e-15*_P23'
.param _P39='1e-14*_P25'
.param _P40='100*_P27'
.param _P41='1e-15*_P29'
.param _P42='1e-14*_P31'
.param _P43='100*_P33'
.param _P44='1e-15*_P35'
.param _P45='V45+V46*radius_+V47*w_'
.param _P46='0.5*(_P45+sqrt(_P45*_P45+0.001))'
.param _P47='V48+V49*radius_+V50*w_'
.param _P48='0.5*(_P47+sqrt(_P47*_P47+0.001))'
.param _P49='100*_P46'
.param _P50='1e-13*_P48'
.param _P51='V51+V52*radius_+V53*w_'
.param _P52='0.5*(_P51+sqrt(_P51*_P51+0.001))'
.param _P53='V54+V55*radius_+V56*w_'
.param _P54='0.5*(_P53+sqrt(_P53*_P53+0.001))'
.param _P55='100*_P52'
.param _P56='1e-13*_P54'
.param _P57='V57+V58*radius_+V59*w_'
.param _P58='0.5*(_P57+sqrt(_P57*_P57+0.001))'
.param _P59='V60+V61*radius_+V62*w_'
.param _P60='0.5*(_P59+sqrt(_P59*_P59+0.001))'
.param _P61='100*_P58'
.param _P62='1e-13*_P60'
cs PLUS MINUS '_P2'
rs1_1 PLUS n1_1 '_P4*(1+drs_2Tdiff_psub)' tc1=0.003
ls1_1 n1_1 ni_1 '_P7*(1+dls_2Tdiff_psub)'
rs2_1 ni_1 n2_1 '_P4*(1+drs_2Tdiff_psub)' tc1=0.003
ls2_1 n2_1 MINUS '_P8*(1+dls_2Tdiff_psub)'
rs1_2 PLUS n1_2 '_P10*(1+drs_2Tdiff_psub)' tc1=0.003
ls1_2 n1_2 MINUS '_P13*(1+dls_2Tdiff_psub)'
k1 ls1_1 ls1_2 K=_P16
k2 ls2_1 ls1_2 K=_P17
c_1_sub PLUS _n1_1_sub '_P36'
rs_1_sub _n1_1_sub PSUB '_P37'
cs_1_sub _n1_1_sub PSUB '_P38'
c_2_sub MINUS _n1_2_sub '_P39'
rs_2_sub _n1_2_sub PSUB '_P40'
cs_2_sub _n1_2_sub PSUB '_P41'
c_3_sub ni_1 _n1_3_sub '_P42'
rs_3_sub _n1_3_sub PSUB '_P43'
cs_3_sub _n1_3_sub PSUB '_P44'
rx_1_2_sub _n1_1_sub _n1_2_sub '_P49'
cx_1_2_sub _n1_1_sub _n1_2_sub '_P50'
rx_1_3_sub _n1_1_sub _n1_3_sub '_P55'
cx_1_3_sub _n1_1_sub _n1_3_sub '_P56'
rx_2_3_sub _n1_2_sub _n1_3_sub '_P61'
cx_2_3_sub _n1_2_sub _n1_3_sub '_P62'
kzero1 ls1_1 ls2_1 K=1e-6
.ends diff_ind_rf_psub
