//* 
//* No part of this file can be released without the consent of SMIC.
//*
//******************************************************************************************
//* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.11
//*
//* Release date       : 4/27/2015
//*
//* Simulation tool    : Cadence Spectre V10.1.1
//*
//*
//*  MOSFET Varactor  :
//*
//*
//*        *--------------------------------------------------------------* 
//*        |                        MOSFET varactor subckt                |     
//*        |==============================================================| 
//*        |   NMOS in NWELL 1.8V      |  pvar18_ckt_rf                   | 
//*        |==============================================================| 
//*        |   NMOS in NWELL 3.3V      |  pvar33_ckt_rf                   | 
//*        *--------------------------------------------------------------*
//*
//*
//*  Junction Diode Varactor  :  
//*
//*        *--------------------------------------------------------------* 
//*        | Junction Diode type   |       1.8V       |        3.3V       |
//*        |==============================================================| 
//*        |       N+/PWELL        |   pvardio18_rf   |   pvardio33_rf    |
//*        *--------------------------------------------------------------*
//*
//*        *--------------------------------------------------------------* 
//*        | Junction Diode subckt |       1.8V       |        3.3V       |
//*        |==============================================================| 
//*        |       N+/PWELL        | pvardio18_ckt_rf | pvardio33_ckt_rf  |
//*        *--------------------------------------------------------------*
//* //*
simulator lang=spectre  insensitive=yes
ahdl_include "gc.va"
//*          
//***************************
//* 0.18um 1.8V MOS Varactor*
//***************************
//* 1=port1, 2=port2
//* Area=Wr*Lr*Nf
subckt pvar18_ckt_rf (1 2)
//* mos varactor scalable model parameters
parameters lr=1u wr=2u nf=12 ar=lr*wr*nf mr=1 mismod_var=1
//* equivalent circuit
+ac0_pvar18_rf     =  0          
+bc0_pvar18_rf     =  3.04e-9    
+cc0_pvar18_rf     =  0  
+geo_var_rf        = ac0_pvar18_rf/(wr*(lr+2.6e-14/lr)*nf*mr)+bc0_pvar18_rf/sqrt(wr*(lr+2.6e-14/lr)*nf*mr)+cc0_pvar18_rf         
+dcgg_pvar18mis_rf = mismod_var*sigma_mis_var_rf*geo_var_rf 
//**subckt parameter              
+rsub1_rf     = max((-629.32*log(nf)+4000), 1e-3) 
+csub1_rf     = max((0.0348*nf+0.1652)*1e-15, 1e-18)
+cox1_rf      = max(((0.004*(lr*1e6)+0.0081)*(wr*1e6)*nf+(0.032*(lr*1e6)+0.0638))*1e-15, 1e-18)
+rsub2_rf     = max((303.64*(lr*1e6)+254.47)*pwr((wr*1e6)*nf,(-0.3054*(lr*1e6)+0.0147)), 1e-3)
+csub2_rf     = max((((0.8728*(lr*1e6)-0.528)*(wr*1e6)+(-3.1644*(lr*1e6)+4.2208))*nf+((-1.7148*(lr*1e6)+4.3055)*(wr*1e6)+(0.6456*(lr*1e6)+1.4517)))*1e-15, 1e-18)
+cox2_rf      = max((((0.126*(lr*1e6)+0.0168)*(wr*1e6)+(0.896*(lr*1e6)+0.828))*nf+((-0.0204*(lr*1e6)+1.4385)*(wr*1e6)+(-0.163*(lr*1e6)+1.0508)))*1e-15, 1e-18)
+djnw_area_rf = (wr*1e6+2*0.12)*(lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*1e-12
+djnw_pj_rf   = (wr*1e6+2*0.12+lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*2*1e-6
+cgg_a2       = a_a2*((8.28*(wr*1e6)*(lr*1e6)*nf+0.4638*(wr*1e6)*nf+0.7149*(lr*1e6)*nf+0.202*(wr*1e6)-0.1569*(lr*1e6)))
+cgg_a1       = a_a1*((1.647*(wr*1e6)*(lr*1e6)*nf+0.4773*(wr*1e6)*nf+0.5422*(lr*1e6)*nf+0.04776*(wr*1e6)+0.01854*(lr*1e6)))
+cgg_x0       = -0.4315*pwr((wr*1e6),-0.07108)*(1-2.758*(lr*1e6)+1.902*(lr*1e6)*(lr*1e6))*pwr(nf+552.3,0.07095*pwr((wr*1e6),0.01743)*pwr((lr*1e6),-1.0097))
+a_a1	      = 1.0704*exp(-0.0385*(lr*1e6))
+a_a2	      = 0.0361*log(lr*1e6)+0.9651
+rs_rf        = max((((((-7.562e-01*(lr*1e6)+1.839e+00)*(wr*1e6)*(wr*1e6)+(6.514e+00*(lr*1e6)-2.316e+01)*(wr*1e6)+(-3.931e+01*(lr*1e6)+1.370e+02))*pwr(nf,((4.100e-03*(lr*1e6)-4.300e-03)*(wr*1e6)*(wr*1e6)+(-4.590e-02*(lr*1e6)+4.900e-02)*(wr*1e6)+(1.446e-01*(lr*1e6)-1.153e+00))))))*(1+drs_pvar18_rf), 1e-6)
//**gate current parameter
+tox    = 1.2518e-08+dtox_pvar18_rf 
+gcie   = 2.449260179                 gcarc = 4.97112503779554                 gcevgc = 1.28405488039671
+gcetc  = 2425.31845182089            gcete = 0.305811750223937                igg_tc = 0.00896             
aigg (22 2) aigg_hdl weff=wr*nf*mr leff=lr+2.6e-14/lr tox=tox gcie=gcie gcarc=gcarc gcevgc=gcevgc gcetc=gcetc gcete=gcete
//* equivalent circuit
ls    (11 22) inductor   l=10p       m=mr    
rs    (1  11) resistor   r=max((((rs_rf*(1+0.04/(v(22,2)*v(22,2)+(0.0004*(wr*1e6)*(wr*1e6)+0.0137*(wr*1e6)+0.4708)*(0.0004*(wr*1e6)*(wr*1e6)+0.0137*(wr*1e6)+0.4708))))*(1+2.266e-03*(temp-25)-3.309e-06*(temp-25)*(temp-25)))), 1e-6) m=mr          
cgg   (22  2) capacitor  c=max((cgg_a2+(cgg_a1-cgg_a2)/(1+exp((v(22,2)-cgg_x0)/((-0.0347*v(22,2)*v(22,2)*v(22,2)*v(22,2)+0.00857*v(22,2)*v(22,2)*v(22,2)+0.131*v(22,2)*v(22,2)-0.0389*v(22,2)+0.19)*(0.00143*(temp-25)+1)))))*(1+dcgg_pvar18_rf)*1e-15, 1e-15) m=mr      
cox1  (1  10) capacitor  c=cox1_rf   m=mr 
rsub1 (10  0) resistor   r=rsub1_rf  m=mr 
csub1 (10  0) capacitor  c=csub1_rf  m=mr 
cox2  (2  20) capacitor  c=cox2_rf   m=mr     
rsub2 (20  0) resistor   r=rsub2_rf  m=mr 
csub2 (20  0) capacitor  c=csub2_rf  m=mr 
djnw  (0   2)
+nwdio_rf
+area  = djnw_area_rf
+pj    = djnw_pj_rf   
+m     = mr      
model nwdio_rf diode
+level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
+dcap = 2 area = 9.6e-009 perim = 4e-004 tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
+is = 2.3733e-006 isw = 2.9142e-014 vb = 15 ibv = 104 
+n = 1.085 ns = 1.085 rs = 8.4602e-009 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
+cj = 0 cjp = 0 vj = 0.41624 vjsw = 0.81575 
+fcs = 0 mj = 0.26295 mjsw = 0.377 fc = 0 
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
+tlev = 1 tlevc = 1 trs = 0.0004 xti = 3 
+cta = 0.0017608 ctp = 0.0012659 pta = 0.00155 ptp = 0.0022128 
+eg = 1.16 
ends pvar18_ckt_rf
//*          
//*************************************
//* 0.18um 3.3V MOS Varactor
//*************************************
//* 1=port1, 2=port2
//* Area=Wr*Lr*Nf
subckt pvar33_ckt_rf (1 2)
//* mos varactor scalable model parameters
parameters lr=1u wr=10u nf=12 ar=lr*wr*nf mr=1 mismod_var=1
//* equivalent circuit
ls    (11 22)  inductor   l=10p
parameters rs_a = (((2.18219600*lr*1e6-1.31073200)*wr*1e6*wr*1e6+(-36.30831000*lr*1e6+23.46962700)*wr*1e6+(106.27523200*lr*1e6-24.91322400))*pwr(nf,((-0.02877400*lr*1e6+0.02830400)*wr*1e6*wr*1e6+(0.40768000*lr*1e6-0.40029000)*wr*1e6+(-1.23126600*lr*1e6+0.17806600))))
parameters rs_b = ((-0.56984200*lr*1e6+0.59987600)*wr*1e6*wr*1e6+(8.46208200*lr*1e6-9.01834500)*wr*1e6+(-27.19727400*lr*1e6+30.22506800))
parameters rs_d = ((-0.05474200*lr*1e6+0.05283200)*wr*1e6*wr*1e6+(0.80293400*lr*1e6-0.77210600)*wr*1e6+(-2.13486200*lr*1e6+2.90342700))
parameters rs_e = ((-0.02549600*lr*1e6+0.03906600)*wr*1e6*wr*1e6+(0.48609400*lr*1e6-0.70076400)*wr*1e6+(-2.59254400*lr*1e6+3.40643400))
// *** mismatch paramters	
+lrr=lr*1e6 wrr=wr*1e6     
+area1 = lrr*wrr*nf        
+geo_var_rf = ac0_pvar33_rf/sqrt(area1*mr)+bc0_pvar33_rf	
+dcgg_pvar33mis_rf = mismod_var*sigma_mis_var_rf*geo_var_rf
rs    (1  11)  resistor   r=max(((rs_a*(1+0.1*rs_e*v(22,2)+0.1*rs_b/(v(22,2)*v(22,2)+rs_d*rs_d)))*(1+2.266E-03*(temp-25)-3.309E-06*(temp-25)*(temp-25)))*(1+drs_pvar33_rf),1e-6) m=mr
rsub1 (10  0)  resistor   r=max((-157.33*log(nf)+1000), 1e-3) m=mr
csub1 (10  0)  capacitor  c=max(((0.058000*lr*1e6+0.131000)*nf+(1.152200*lr*1e6+0.263900))*1e-15, 1e-18) m=mr
cox1  (1  10)  capacitor  c=max((((-0.02130818*lr*1e6+0.02299185)*wr*1e6+(0.19167958*lr*1e6-0.03172040))*nf+(-0.01930408*lr*1e6+0.02256428)*wr*1e6+(0.03578980*lr*1e6-0.12376429))*1e-15, 1e-18) m=mr
rsub2 (20  0)  resistor   r=max(((0.17509600*lr*1e6+0.13622500)*wr*1e6+(-3.13181000*lr*1e6-5.98751100))*nf+(-0.36204000*lr*1e6-16.93326600)*wr*1e6+(-5.25510200*lr*1e6+ 419.97183700), 1e-3) m=mr
csub2 (20  0)  capacitor  c=max((((-0.05913800*lr*1e6+3.56503100)*wr*1e6+(2.06525200*lr*1e6+0.32525500))*pwr(nf,((0.02163000*lr*1e6-0.05084700)*wr*1e6+(-0.18202800*lr*1e6+0.69376000))))*1e-15, 1e-18) m=mr
cox2  (2  20)  capacitor  c=max((((0.03803200*lr*1e6+0.07406700)*wr*1e6+(1.19708000*lr*1e6+0.60749200))*nf+(0.10622800*lr*1e6+1.37163800)*wr*1e6+(-0.25722800*lr*1e6+1.02081900))*1e-15, 1e-18) m=mr
djnw (0    2) nwdio_rf area=(wr*1e6+2*0.12)*(lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*1e-12  pj=(wr*1e6+2*0.12+lr*1e6*nf+(nf-1)*0.54+2*0.48+2*0.12)*2*1e-6 m=mr
parameters cgg_a1     = a_a1*((4.924416e+00*lr*1e6+3.885705e-01)*wr*1e6*nf+(5.756613e-02*lr*1e6+3.680246e-01))
parameters cgg_a2     = a_a2*((1.490944e+00*lr*1e6+4.324138e-01)*wr*1e6*nf+(-9.410417e-02*lr*1e6+3.779284e-01))
parameters cgg_x0     = (-(-2.510018e-02*lr*1e6+2.329891e-01)*pwr(wr*1e6*nf,(2.091532e-02*lr*1e6-2.966834e-02)))
parameters cgg_dx     = (-(3.454607e-02*lr*1e6+3.079878e-01)*pwr(wr*1e6*nf,(-1.125777e-02*lr*1e6+2.882598e-03)))
parameters a_a1	= (1.0147*pwr(wr*1e6,-0.0211))
parameters a_a2	= (1.0+0.0157*log(nf))
cgg   (22  2)  capacitor  c=max(((cgg_a2+(cgg_a1-cgg_a2)/(1+exp((v(22,2)-cgg_x0)/(cgg_dx*(0.00143*(temp-25)+1))))))*(1+dcgg_pvar33mis_rf)*(1+dcgg_pvar33_rf)*1e-15, 1e-15) m=mr
//model nwdio_rf diode
//+level = 1 is = 1.42e-06 allow_scaling = yes dskip = no imax=1e20 isw = 1.00e-15 
//+n = 1.0128 ns = 1.0128 rs = 2.44e-08 ik = 1.1e+04 ikp = 7.75e-06 
//+bv = 15.0 ibv = 104.2 
//+trs = 9.47e-04 eg = 1.16 tnom = 25.0 
//+xti = 3.0 cjo = 0 mj = 0.317 
//+vj = 0.494 cjsw = 0 mjsw = 0.383 
//+vjsw = 0.9 cta = 0.002 ctp = 0.00121 
//+pta = 0.00253 ptp = 0.00217 tlev = 1 
//+tlevc = 1
//+fc = 0 
model nwdio_rf diode
parameters level = 1 allow_scaling = yes dskip = no imax = 1e20  minr = 1e-6
// **************************************************************
// *               GENERAL PARAMETERS
// **************************************************************
parameters dcap = 2 area = 9.6e-009 perim = 4e-004
// tnom = 25 
// **************************************************************
// *               DC PARAMETERS
// **************************************************************
parameters is = 2.3733e-006 isw = 2.9142e-014 vb = 15 ibv = 104 
parameters n = 1.085 ns = 1.085 rs = 8.4602e-009 
// **************************************************************
// *               CAPACITANCE PARAMETERS
// **************************************************************
parameters cj = 0 cjp = 0 vj = 0.41624 vjsw = 0.81575 
parameters fcs = 0 mj = 0.26295 mjsw = 0.377 fc = 0 
// **************************************************************
// *               NOISE PARAMETERS
// **************************************************************
// **************************************************************
// *               TEMPERATURE PARAMETERS
// **************************************************************
parameters tlev = 1 tlevc = 1 trs = 0.0004 xti = 3 
parameters cta = 0.0017608 ctp = 0.0012659 pta = 0.00155 ptp = 0.0022128 
parameters eg = 1.16 
ends pvar33_ckt_rf
//*
//****************************
//* 0.18um 1.8V P+/NW Varactor
//****************************
//* 1=port1, 2=port2
//* Area=Wr*Lr*Nf
subckt pvardio18_ckt_rf (1 2)
//* P+/NW junction varactor scalable model parameters
parameters lr=20u wr=5u nf=10 ar=lr*wr*nf pj=(lr+wr)*2*nf
//* equivalent circuit
ls    (1 11)  inductor   l=(0.07947+(1.7134E-05*ar*1E12)-(3.865E-09*ar*ar*1E24))*1E-9       
rs    (11 22) resistor   r=0.23268+(3.334E+03/(ar*1E12))+(8.9147E+04/(ar*ar*1E24))
rsub1 (10 0)  resistor   r=1E+05
csub1 (10 0)  capacitor  c=1*1E-15
cox1  (1 10)  capacitor  c=1*1E-15  
rsub2 (20 0)  resistor   r=1940-(1.6342*ar*1E12)+(4.2816E-04*ar*ar*1E24)
csub2 (20 0)  capacitor  c=(2.75025+(2.787E-03*ar*1E12)+(1.3682E-06*ar*ar*1E24))*1E-15        
cox2  (2 20)  capacitor  c=(27.96263+(0.53519*ar*1E12)-(9.0589E-05*ar*ar*1E24))*1E-15
diode (22 2)  pvardio18_rf area=ar pj=pj
//* P+/Nwell varactor model
model pvardio18_rf diode
+level = 1 is = 1.1913E-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15
+cjo = 1.1495e-3 mj = 0.37316 
+tnom = 25 vj = 0.76958 cta = 0.000876 
+pta = 0.00153 fc = 0 
+eg = 1.16 tlev = 1 tlevc = 1
+n = 0.98812 ns = 0.98812 rs = 0 ik = 4.2216e+06 ikp = 2.43E-03 
+bv = 12 ibv = 2000 trs = 1.78e-03  xti = 3.0 
ends pvardio18_ckt_rf
//*
//****************************
//* 0.18um 3.3V P+/NW Varactor
//****************************
//* 1=port1, 2=port2
//* Area=Wr*Lr*Nf
subckt pvardio33_ckt_rf (1 2)
//* P+/NW junction varactor scalable model parameters
parameters lr=20u wr=5u nf=10 ar=lr*wr*nf  pj=(lr+wr)*2*nf
//* equivalent circuit
ls    (1 11)  inductor   l=(0.08203+(1.3302E-05*ar*1E12)-(1.844E-09*ar*ar*1E24))*1E-9       
rs    (11 22) resistor   r=0.25902+(3.3475E+03/(ar*1E12))+(1.0295E+05/(ar*ar*1E24))
rsub1 (10 0)  resistor   r=1E+05
csub1 (10 0)  capacitor  c=1*1E-15
cox1  (1 10)  capacitor  c=1*1E-15  
rsub2 (20 0)  resistor   r=1.869E+03-(1.49373*ar*1E12)+(3.7877E-04*ar*ar*1E24)
csub2 (20 0)  capacitor  c=(3.81691-(1.5322E-03*ar*1E12)+(4.0789E-06*ar*ar*1E24))*1E-15        
cox2  (2 20)  capacitor  c=(64.90675+(0.37036*ar*1E12)+(1.0985E-06*ar*ar*1E24))*1E-15
diode (22 2)  pvardio33_rf area=ar pj=pj
//* P+/Nwell varactor model
model pvardio33_rf diode
+level = 1 is = 1.3141E-07 allow_scaling = yes dskip = no imax=1e20 isw = 1e-15
+cjo = 1.1455E-3  mj = 0.3793 
+tnom = 25 vj = 0.792 cta = 0.000897
+pta = 0.00166 fc = 0 
+eg = 1.16 tlev = 1 tlevc = 1 
+n = 0.99195 ns = 0.99195 rs = 0 ik = 4.5171E+06  
+bv = 12 ibv = 2000 xti = 3.0  trs = 1.24e-03 ikp = 2.42e-03
ends pvardio33_ckt_rf
//*
